
module HFC1 (N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670, N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873);

input N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670;
output N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873;
  wire   N1118, N226, N935, N1282, N1142, N1511, N1401, N258, N733, N1479,
         N1330, N423, N2, N77, N124, N227, N249, N287, N416, N513, N528, N678,
         N684, N749, N882, N949, N1074, N1091, N1104, N1134, N1136, N1273,
         N1332, N1405, N1502, N1670, N264, N1012, N383, N1221, N736, N8, N191,
         N1549, N911, N1246, N1513, N1117, N422, N1293, N93, N751, N1123,
         N1077, N142, N389, N1131, N1115, N544, N1406, N510, N1773, N562,
         N1664, N1711, N254, N1362, N1331, N762, N174, N938, N235, N841, N660,
         N67, N954, N520, N1766, N1138, N1869, N811, N330, N884, N1812, N823,
         N1522, N166, N1259, N984, N740, N1786, N501, N31, N1011, N344, N1756,
         N722, N63, N1596, N1066, N304, N800, N979, N150, N550, N534, N1605,
         N1477, N1297, N425, N1587, N502, N1161, N1010, N628, N1651, N35, N117,
         N59, N402, N1346, N605, N414, N1544, N1452, N1408, N1636, N750, N1767,
         N1491, N1127, N673, N52, N1232, N1483, N1385, N1277, N1485, N1496,
         N621, N1714, N1063, N1447, N1826, N1300, N487, N365, N24, N1838,
         N1823, N102, N230, N824, N408, N1113, N1600, N1099, N1047, N707,
         N1410, N873, N79, N234, N897, N744, N1309, N955, N1359, N732, N74,
         N781, N647, N1050, N292, N242, N922, N1320, N598, N1634, N1165, N1561,
         N685, N38, N617, N1722, N1662, N42, N1667, N1685, N623, N1159, N1205,
         N1648, N1235, N1179, N294, N229, N1768, N288, N1602, N223, N1214,
         N724, N925, N1507, N972, N415, N939, N1218, N1239, N1687, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435;
  assign N847 = N1118;
  assign N237 = N226;
  assign N735 = N935;
  assign N1046 = N1282;
  assign N940 = N1142;
  assign N361 = N1511;
  assign N1769 = N1401;
  assign N1497 = N1401;
  assign N1265 = N1401;
  assign N928 = N1401;
  assign N209 = N1401;
  assign N347 = N1401;
  assign N585 = N1401;
  assign N729 = N1401;
  assign N825 = N258;
  assign N891 = N733;
  assign N348 = N733;
  assign N1069 = N733;
  assign N675 = N733;
  assign N381 = N1479;
  assign N350 = N1330;
  assign N1445 = N423;
  assign N357 = N423;
  assign N316 = N423;
  assign N377 = N423;
  assign N871 = N2;
  assign N1870 = N2;
  assign N946 = N2;
  assign N569 = N2;
  assign N860 = N77;
  assign N181 = N124;
  assign N1772 = N124;
  assign N761 = N124;
  assign N110 = N124;
  assign N163 = N227;
  assign N1465 = N227;
  assign N1286 = N227;
  assign N721 = N227;
  assign N780 = N249;
  assign N1841 = N249;
  assign N1347 = N249;
  assign N1310 = N249;
  assign N111 = N249;
  assign N980 = N287;
  assign N584 = N287;
  assign N413 = N287;
  assign N14 = N287;
  assign N252 = N416;
  assign N794 = N416;
  assign N481 = N416;
  assign N431 = N416;
  assign N275 = N416;
  assign N274 = N513;
  assign N1489 = N513;
  assign N1440 = N513;
  assign N107 = N513;
  assign N387 = N528;
  assign N1125 = N528;
  assign N801 = N528;
  assign N509 = N528;
  assign N1822 = N678;
  assign N1379 = N678;
  assign N664 = N684;
  assign N1444 = N684;
  assign N1255 = N684;
  assign N392 = N684;
  assign N167 = N684;
  assign N495 = N749;
  assign N403 = N749;
  assign N1438 = N882;
  assign N18 = N882;
  assign N43 = N949;
  assign N39 = N949;
  assign N1640 = N1074;
  assign N1560 = N1074;
  assign N1471 = N1074;
  assign N1013 = N1074;
  assign N1606 = N1091;
  assign N1791 = N1091;
  assign N1001 = N1091;
  assign N478 = N1091;
  assign N368 = N1091;
  assign N217 = N1091;
  assign N1071 = N1104;
  assign N633 = N1104;
  assign N69 = N1104;
  assign N5 = N1104;
  assign N1325 = N1134;
  assign N839 = N1134;
  assign N869 = N1136;
  assign N1552 = N1136;
  assign N1433 = N1136;
  assign N1350 = N1136;
  assign N952 = N1136;
  assign N1547 = N1273;
  assign N1197 = N1273;
  assign N91 = N1332;
  assign N1720 = N1332;
  assign N1256 = N1332;
  assign N1110 = N1332;
  assign N642 = N1332;
  assign N358 = N1332;
  assign N1199 = N1405;
  assign N1675 = N1405;
  assign N687 = N1405;
  assign N57 = N1405;
  assign N1737 = N1502;
  assign N1594 = N1502;
  assign N136 = N1502;
  assign N1775 = N1670;
  assign N1514 = N1670;
  assign N1075 = N1670;
  assign N272 = N1670;
  assign N83 = N1670;
  assign N1859 = N264;
  assign N137 = N264;
  assign N1170 = N1012;
  assign N680 = N1012;
  assign N681 = N383;
  assign N615 = N383;
  assign N251 = N383;
  assign N821 = N383;
  assign N1194 = N1221;
  assign N921 = N1221;
  assign N1508 = N736;
  assign N106 = N8;
  assign N1842 = N191;
  assign N1450 = N1549;
  assign N165 = N1549;
  assign N177 = N911;
  assign N1240 = N1246;
  assign N333 = N1513;
  assign N1659 = N1117;
  assign N1067 = N1117;
  assign N899 = N422;
  assign N1789 = N1293;
  assign N894 = N1293;
  assign N1383 = N93;
  assign N1400 = N751;
  assign N1052 = N751;
  assign N445 = N751;
  assign N1089 = N751;
  assign N620 = N751;
  assign N1421 = N1123;
  assign N1654 = N1077;
  assign N1749 = N142;
  assign N1112 = N142;
  assign N281 = N142;
  assign N190 = N142;
  assign N178 = N142;
  assign N1301 = N389;
  assign N1076 = N389;
  assign N926 = N389;
  assign N629 = N389;
  assign N1079 = N389;
  assign N1480 = N1131;
  assign N1467 = N1115;
  assign N782 = N544;
  assign N1436 = N1406;
  assign N1343 = N1406;
  assign N374 = N1406;
  assign N816 = N1406;
  assign N10 = N1406;
  assign N1620 = N510;
  assign N218 = N510;
  assign N1472 = N1773;
  assign N1751 = N562;
  assign N1361 = N562;
  assign N656 = N562;
  assign N22 = N562;
  assign N554 = N562;
  assign N1840 = N1664;
  assign N1060 = N1664;
  assign N1716 = N1711;
  assign N1404 = N1711;
  assign N151 = N1711;
  assign N314 = N1711;
  assign N655 = N1711;
  assign N969 = N1711;
  assign N1323 = N254;
  assign N852 = N254;
  assign N557 = N254;
  assign N428 = N254;
  assign N188 = N254;
  assign N1683 = N254;
  assign N1002 = N1362;
  assign N12 = N1362;
  assign N1671 = N1331;
  assign N1177 = N1331;
  assign N679 = N1331;
  assign N33 = N1331;
  assign N1416 = N1331;
  assign N779 = N762;
  assign N483 = N174;
  assign N100 = N174;
  assign N335 = N938;
  assign N959 = N938;
  assign N1295 = N235;
  assign N323 = N841;
  assign N220 = N841;
  assign N94 = N841;
  assign N80 = N841;
  assign N26 = N841;
  assign N1032 = N841;
  assign N1145 = N841;
  assign N683 = N841;
  assign N688 = N841;
  assign N433 = N660;
  assign N1643 = N67;
  assign N1595 = N67;
  assign N690 = N67;
  assign N211 = N67;
  assign N109 = N67;
  assign N311 = N67;
  assign N1843 = N954;
  assign N1808 = N520;
  assign N1752 = N520;
  assign N1478 = N520;
  assign N505 = N520;
  assign N202 = N520;
  assign N401 = N1766;
  assign N1754 = N1138;
  assign N1186 = N1138;
  assign N391 = N1138;
  assign N135 = N1138;
  assign N981 = N1138;
  assign N822 = N1869;
  assign N596 = N1869;
  assign N1863 = N811;
  assign N1741 = N811;
  assign N1412 = N811;
  assign N815 = N811;
  assign N315 = N811;
  assign N337 = N811;
  assign N1796 = N330;
  assign N1014 = N330;
  assign N1619 = N884;
  assign N1833 = N884;
  assign N320 = N1812;
  assign N50 = N1812;
  assign N1469 = N823;
  assign N1614 = N1522;
  assign N1085 = N1522;
  assign N1162 = N166;
  assign N798 = N166;
  assign N419 = N1259;
  assign N1088 = N1259;
  assign N970 = N984;
  assign N295 = N984;
  assign N121 = N984;
  assign N1409 = N984;
  assign N1128 = N740;
  assign N1003 = N740;
  assign N988 = N740;
  assign N958 = N740;
  assign N720 = N740;
  assign N438 = N740;
  assign N1627 = N740;
  assign N583 = N1786;
  assign N169 = N1786;
  assign N1686 = N501;
  assign N1395 = N501;
  assign N1538 = N31;
  assign N1023 = N31;
  assign N831 = N31;
  assign N1036 = N31;
  assign N775 = N1011;
  assign N65 = N1011;
  assign N1798 = N344;
  assign N1617 = N344;
  assign N407 = N1756;
  assign N944 = N722;
  assign N723 = N63;
  assign N1858 = N1596;
  assign N696 = N1596;
  assign N631 = N1596;
  assign N577 = N1596;
  assign N1718 = N1596;
  assign N1555 = N1066;
  assign N658 = N1066;
  assign N1490 = N304;
  assign N1846 = N800;
  assign N1811 = N800;
  assign N1689 = N800;
  assign N1238 = N800;
  assign N1193 = N800;
  assign N697 = N800;
  assign N7 = N800;
  assign N1747 = N800;
  assign N1082 = N979;
  assign N659 = N979;
  assign N340 = N979;
  assign N973 = N979;
  assign N1120 = N150;
  assign N1098 = N150;
  assign N158 = N150;
  assign N1607 = N550;
  assign N931 = N534;
  assign N498 = N534;
  assign N471 = N534;
  assign N173 = N534;
  assign N30 = N534;
  assign N1169 = N534;
  assign N253 = N1605;
  assign N1303 = N1477;
  assign N974 = N1297;
  assign N1080 = N425;
  assign N634 = N1587;
  assign N40 = N502;
  assign N1463 = N1161;
  assign N1777 = N1010;
  assign N260 = N628;
  assign N613 = N1651;
  assign N758 = N35;
  assign N573 = N117;
  assign N1785 = N59;
  assign N430 = N402;
  assign N224 = N1346;
  assign N1377 = N605;
  assign N159 = N414;
  assign N565 = N414;
  assign N360 = N1544;
  assign N160 = N1452;
  assign N1744 = N1408;
  assign N1188 = N1636;
  assign N1418 = N750;
  assign N1364 = N1767;
  assign N469 = N1767;
  assign N746 = N1491;
  assign N813 = N1127;
  assign N1215 = N673;
  assign N305 = N52;
  assign N319 = N1232;
  assign N266 = N1483;
  assign N759 = N1385;
  assign N436 = N1277;
  assign N129 = N1485;
  assign N298 = N1496;
  assign N1787 = N621;
  assign N406 = N1714;
  assign N699 = N1063;
  assign N228 = N1447;
  assign N32 = N1826;
  assign N592 = N1300;
  assign N1318 = N1300;
  assign N622 = N1300;
  assign N132 = N487;
  assign N157 = N365;
  assign N561 = N24;
  assign N769 = N1838;
  assign N1526 = N1823;
  assign N1696 = N102;
  assign N662 = N230;
  assign N309 = N824;
  assign N301 = N824;
  assign N246 = N408;
  assign N1609 = N1113;
  assign N250 = N1113;
  assign N819 = N1600;
  assign N555 = N1099;
  assign N1027 = N1047;
  assign N105 = N1047;
  assign N189 = N707;
  assign N1093 = N1410;
  assign N396 = N1410;
  assign N1518 = N873;
  assign N21 = N79;
  assign N1183 = N234;
  assign N1064 = N897;
  assign N1029 = N744;
  assign N540 = N744;
  assign N950 = N1309;
  assign N162 = N1309;
  assign N421 = N955;
  assign N96 = N955;
  assign N1389 = N1359;
  assign N1070 = N1359;
  assign N1005 = N1359;
  assign N473 = N1359;
  assign N336 = N1359;
  assign N270 = N732;
  assign N334 = N74;
  assign N1430 = N781;
  assign N204 = N647;
  assign N1153 = N1050;
  assign N200 = N292;
  assign N1353 = N292;
  assign N1503 = N242;
  assign N808 = N922;
  assign N90 = N1320;
  assign N104 = N1320;
  assign N892 = N598;
  assign N1210 = N1634;
  assign N576 = N1165;
  assign N331 = N1561;
  assign N1509 = N685;
  assign N1229 = N38;
  assign N497 = N617;
  assign N551 = N1722;
  assign N1216 = N1662;
  assign N625 = N42;
  assign N1155 = N1667;
  assign N247 = N1685;
  assign N1236 = N623;
  assign N297 = N1159;
  assign N682 = N1205;
  assign N168 = N1648;
  assign N861 = N1235;
  assign N199 = N1179;
  assign N1545 = N294;
  assign N134 = N229;
  assign N455 = N1768;
  assign N885 = N288;
  assign N302 = N288;
  assign N1571 = N288;
  assign N1825 = N1602;
  assign N703 = N1602;
  assign N739 = N223;
  assign N370 = N223;
  assign N1037 = N1214;
  assign N708 = N1214;
  assign N98 = N724;
  assign N16 = N724;
  assign N122 = N925;
  assign N803 = N1507;
  assign N1810 = N1507;
  assign N1103 = N972;
  assign N214 = N415;
  assign N193 = N939;
  assign N255 = N1218;
  assign N717 = N1239;
  assign N627 = N1687;

  CKND2D0BWPHVT U470 ( .A1(N310), .A2(N383), .ZN(N987) );
  CKND2D0BWPHVT U471 ( .A1(N783), .A2(N1331), .ZN(N95) );
  AN2D0BWPHVT U472 ( .A1(N142), .A2(N171), .Z(N934) );
  CKND2D0BWPHVT U473 ( .A1(N954), .A2(N389), .ZN(N897) );
  CKND2D0BWPHVT U474 ( .A1(N1800), .A2(N287), .ZN(N858) );
  CKND2D0BWPHVT U475 ( .A1(N951), .A2(N435), .ZN(N82) );
  CKND2D0BWPHVT U476 ( .A1(N179), .A2(N1331), .ZN(N951) );
  CKND2D0BWPHVT U477 ( .A1(N1015), .A2(N1596), .ZN(N796) );
  CKND2D0BWPHVT U478 ( .A1(N884), .A2(N1237), .ZN(N787) );
  CKND2D0BWPHVT U479 ( .A1(N1767), .A2(N1507), .ZN(N750) );
  CKND2D0BWPHVT U480 ( .A1(N865), .A2(N1138), .ZN(N68) );
  CKND2D0BWPHVT U481 ( .A1(N206), .A2(N416), .ZN(N667) );
  CKND2D0BWPHVT U482 ( .A1(N991), .A2(N1000), .ZN(N657) );
  CKND2D0BWPHVT U483 ( .A1(N59), .A2(N227), .ZN(N991) );
  CKND2D0BWPHVT U484 ( .A1(N1479), .A2(N568), .ZN(N651) );
  CKND2D0BWPHVT U485 ( .A1(N249), .A2(N1011), .ZN(N647) );
  AN2D0BWPHVT U486 ( .A1(N142), .A2(N578), .Z(N635) );
  CKND2D0BWPHVT U487 ( .A1(N984), .A2(N626), .ZN(N62) );
  CKND2D0BWPHVT U488 ( .A1(N1722), .A2(N1670), .ZN(N617) );
  CKND2D0BWPHVT U489 ( .A1(N235), .A2(N1259), .ZN(N598) );
  CKND2D0BWPHVT U490 ( .A1(N994), .A2(N1357), .ZN(N578) );
  CKND2D0BWPHVT U491 ( .A1(N590), .A2(N914), .ZN(N994) );
  CKND0BWPHVT U492 ( .I(N804), .ZN(N914) );
  CKND0BWPHVT U493 ( .I(N1179), .ZN(N590) );
  CKND2D0BWPHVT U494 ( .A1(N859), .A2(N1092), .ZN(N538) );
  CKND2D0BWPHVT U495 ( .A1(N117), .A2(N124), .ZN(N859) );
  CKND2D0BWPHVT U496 ( .A1(N1786), .A2(N1664), .ZN(N500) );
  CKND2D0BWPHVT U497 ( .A1(N744), .A2(N288), .ZN(N494) );
  CKND2D0BWPHVT U498 ( .A1(N870), .A2(N1136), .ZN(N447) );
  CKND2D0BWPHVT U499 ( .A1(N810), .A2(N2), .ZN(N439) );
  CKND2D0BWPHVT U500 ( .A1(N35), .A2(N287), .ZN(N435) );
  CKND2D0BWPHVT U501 ( .A1(N660), .A2(N534), .ZN(N38) );
  CKND0BWPHVT U502 ( .I(N546), .ZN(N364) );
  CKND2D0BWPHVT U503 ( .A1(N964), .A2(N948), .ZN(N363) );
  CKND2D0BWPHVT U504 ( .A1(N300), .A2(N1138), .ZN(N948) );
  CKND2D0BWPHVT U505 ( .A1(N425), .A2(N528), .ZN(N964) );
  AN2D0BWPHVT U506 ( .A1(N142), .A2(N616), .Z(N325) );
  CKND2D0BWPHVT U507 ( .A1(N900), .A2(N1264), .ZN(N616) );
  CKND2D0BWPHVT U508 ( .A1(N422), .A2(N645), .ZN(N900) );
  CKND0BWPHVT U509 ( .I(N1623), .ZN(N645) );
  CKND0BWPHVT U510 ( .I(N226), .ZN(N422) );
  CKND2D0BWPHVT U511 ( .A1(N593), .A2(N349), .ZN(N313) );
  CKND2D0BWPHVT U512 ( .A1(N1474), .A2(N1780), .ZN(N349) );
  CKND2D0BWPHVT U513 ( .A1(N726), .A2(N1033), .ZN(N593) );
  CKND2D0BWPHVT U514 ( .A1(N609), .A2(N296), .ZN(N307) );
  CKND2D0BWPHVT U515 ( .A1(N1763), .A2(N254), .ZN(N609) );
  CKND2D0BWPHVT U516 ( .A1(N1161), .A2(N249), .ZN(N296) );
  CKND2D0BWPHVT U517 ( .A1(N1786), .A2(N811), .ZN(N294) );
  CKND2D0BWPHVT U518 ( .A1(N486), .A2(N528), .ZN(N265) );
  CKND2D0BWPHVT U519 ( .A1(N1667), .A2(N124), .ZN(N230) );
  CKND2D0BWPHVT U520 ( .A1(N542), .A2(N1151), .ZN(N221) );
  CKND2D0BWPHVT U521 ( .A1(N933), .A2(N800), .ZN(N542) );
  CKND2D0BWPHVT U522 ( .A1(N641), .A2(N282), .ZN(N1850) );
  CKND2D0BWPHVT U523 ( .A1(N1202), .A2(N534), .ZN(N282) );
  CKND2D0BWPHVT U524 ( .A1(N1477), .A2(N1670), .ZN(N641) );
  CKND0BWPHVT U525 ( .I(N288), .ZN(N1786) );
  CKND2D0BWPHVT U526 ( .A1(N824), .A2(N1742), .ZN(N1781) );
  CKND0BWPHVT U527 ( .I(N726), .ZN(N1780) );
  CKND2D0BWPHVT U528 ( .A1(N1417), .A2(N1502), .ZN(N726) );
  CKND2D0BWPHVT U529 ( .A1(N908), .A2(N343), .ZN(N171) );
  CKND2D0BWPHVT U530 ( .A1(N400), .A2(N234), .ZN(N343) );
  CKND2D0BWPHVT U531 ( .A1(N1799), .A2(N354), .ZN(N908) );
  CKND0BWPHVT U532 ( .I(N400), .ZN(N354) );
  CKND2D0BWPHVT U533 ( .A1(n419), .A2(N949), .ZN(N400) );
  CKND0BWPHVT U534 ( .I(N234), .ZN(N1799) );
  CKND2D0BWPHVT U535 ( .A1(N649), .A2(N604), .ZN(N1681) );
  CKND2D0BWPHVT U536 ( .A1(N728), .A2(N811), .ZN(N604) );
  CKND2D0BWPHVT U537 ( .A1(N1346), .A2(N684), .ZN(N649) );
  CKND2D0BWPHVT U538 ( .A1(N1266), .A2(N544), .ZN(N1669) );
  CKND2D0BWPHVT U539 ( .A1(N722), .A2(N911), .ZN(N1636) );
  CKND0BWPHVT U540 ( .I(N1507), .ZN(N722) );
  CKND2D0BWPHVT U541 ( .A1(N1768), .A2(N1165), .ZN(N1634) );
  CKND2D0BWPHVT U542 ( .A1(N814), .A2(N128), .ZN(N1506) );
  CKND2D0BWPHVT U543 ( .A1(N1651), .A2(N1405), .ZN(N814) );
  CKND2D0BWPHVT U544 ( .A1(N1123), .A2(N254), .ZN(N1496) );
  CKND2D0BWPHVT U545 ( .A1(N621), .A2(N249), .ZN(N1485) );
  AN2D0BWPHVT U546 ( .A1(N142), .A2(N589), .Z(N1484) );
  CKND2D0BWPHVT U547 ( .A1(N437), .A2(N388), .ZN(N589) );
  CKND2D0BWPHVT U548 ( .A1(N492), .A2(N1362), .ZN(N388) );
  CKND2D0BWPHVT U549 ( .A1(N258), .A2(N356), .ZN(N437) );
  CKND0BWPHVT U550 ( .I(N492), .ZN(N356) );
  XNR2D0BWPHVT U551 ( .A1(N1266), .A2(N824), .ZN(N492) );
  CKND0BWPHVT U552 ( .I(N1033), .ZN(N1474) );
  CKND2D0BWPHVT U553 ( .A1(N1288), .A2(N1268), .ZN(N1448) );
  CKND2D0BWPHVT U554 ( .A1(N874), .A2(N1499), .ZN(N1424) );
  CKND2D0BWPHVT U555 ( .A1(N1587), .A2(N416), .ZN(N1499) );
  CKND2D0BWPHVT U556 ( .A1(N1152), .A2(N67), .ZN(N874) );
  NR2D0BWPHVT U557 ( .A1(N523), .A2(N1342), .ZN(N1423) );
  AN4D0BWPHVT U558 ( .A1(N827), .A2(N248), .A3(N77), .A4(N150), .Z(N523) );
  INR2D0BWPHVT U559 ( .A1(N1563), .B1(N1283), .ZN(N827) );
  AN4D0BWPHVT U560 ( .A1(N1158), .A2(N1190), .A3(n420), .A4(n421), .Z(N1563)
         );
  AN4D0BWPHVT U561 ( .A1(N380), .A2(N318), .A3(N1736), .A4(N1532), .Z(n421) );
  ND3D0BWPHVT U562 ( .A1(N1146), .A2(N1501), .A3(n422), .ZN(N1532) );
  ND3D0BWPHVT U563 ( .A1(N341), .A2(N1429), .A3(n422), .ZN(N1736) );
  ND3D0BWPHVT U564 ( .A1(n423), .A2(N630), .A3(N61), .ZN(N318) );
  NR2D0BWPHVT U565 ( .A1(N1063), .A2(N781), .ZN(N61) );
  ND3D0BWPHVT U566 ( .A1(N630), .A2(N264), .A3(n423), .ZN(N380) );
  AN2D0BWPHVT U567 ( .A1(N1494), .A2(N1326), .Z(n420) );
  ND3D0BWPHVT U568 ( .A1(N1757), .A2(N1501), .A3(n422), .ZN(N1494) );
  AN2D0BWPHVT U569 ( .A1(N142), .A2(N993), .Z(N1419) );
  CKND2D0BWPHVT U570 ( .A1(N379), .A2(N1562), .ZN(N993) );
  CKND2D0BWPHVT U571 ( .A1(N971), .A2(N1408), .ZN(N1562) );
  CKND2D0BWPHVT U572 ( .A1(N278), .A2(N663), .ZN(N379) );
  CKND0BWPHVT U573 ( .I(N971), .ZN(N663) );
  CKND2D0BWPHVT U574 ( .A1(n419), .A2(N678), .ZN(N971) );
  CKND0BWPHVT U575 ( .I(N1408), .ZN(N278) );
  CKND2D0BWPHVT U576 ( .A1(N1053), .A2(N1048), .ZN(N1417) );
  CKND2D0BWPHVT U577 ( .A1(N97), .A2(N595), .ZN(N1358) );
  CKND2D0BWPHVT U578 ( .A1(N1388), .A2(N180), .ZN(N595) );
  CKND0BWPHVT U579 ( .I(N212), .ZN(N180) );
  CKND0BWPHVT U580 ( .I(N19), .ZN(N1388) );
  CKND2D0BWPHVT U581 ( .A1(N212), .A2(N19), .ZN(N97) );
  CKND2D0BWPHVT U582 ( .A1(N842), .A2(N1398), .ZN(N19) );
  CKND2D0BWPHVT U583 ( .A1(N531), .A2(N1333), .ZN(N1398) );
  CKND0BWPHVT U584 ( .I(N1025), .ZN(N531) );
  CKND2D0BWPHVT U585 ( .A1(N1676), .A2(N1025), .ZN(N842) );
  CKND0BWPHVT U586 ( .I(N1333), .ZN(N1676) );
  CKND2D0BWPHVT U587 ( .A1(N953), .A2(N1502), .ZN(N212) );
  CKND2D0BWPHVT U588 ( .A1(N1141), .A2(N904), .ZN(N953) );
  CKND2D0BWPHVT U589 ( .A1(N804), .A2(N1179), .ZN(N1357) );
  CKND2D0BWPHVT U590 ( .A1(n419), .A2(N174), .ZN(N804) );
  INR3D0BWPHVT U591 ( .A1(N248), .B1(N1502), .B2(N77), .ZN(N1342) );
  ND4D0BWPHVT U592 ( .A1(N326), .A2(N1501), .A3(N1429), .A4(N630), .ZN(N248)
         );
  CKND2D0BWPHVT U593 ( .A1(N546), .A2(N519), .ZN(N1333) );
  XNR2D0BWPHVT U594 ( .A1(N1664), .A2(N288), .ZN(N546) );
  ND3D0BWPHVT U595 ( .A1(N72), .A2(N1429), .A3(n422), .ZN(N1326) );
  AN3D0BWPHVT U596 ( .A1(N630), .A2(N131), .A3(N326), .Z(n422) );
  CKND2D0BWPHVT U597 ( .A1(N938), .A2(N1300), .ZN(N1298) );
  CKND2D0BWPHVT U598 ( .A1(N909), .A2(N984), .ZN(N1288) );
  CKND2D0BWPHVT U599 ( .A1(N743), .A2(N979), .ZN(N128) );
  CKND2D0BWPHVT U600 ( .A1(N284), .A2(N125), .ZN(N1279) );
  CKND2D0BWPHVT U601 ( .A1(N712), .A2(N520), .ZN(N284) );
  CKND2D0BWPHVT U602 ( .A1(N628), .A2(N1074), .ZN(N1268) );
  CKND0BWPHVT U603 ( .I(N1742), .ZN(N1266) );
  CKND2D0BWPHVT U604 ( .A1(n419), .A2(N882), .ZN(N1742) );
  CKND2D0BWPHVT U605 ( .A1(N1623), .A2(N226), .ZN(N1264) );
  CKND2D0BWPHVT U606 ( .A1(n419), .A2(N344), .ZN(N1623) );
  CKND0BWPHVT U607 ( .I(N1768), .ZN(N1259) );
  CKND2D0BWPHVT U608 ( .A1(N1297), .A2(N513), .ZN(N125) );
  CKND2D0BWPHVT U609 ( .A1(N288), .A2(N684), .ZN(N1235) );
  CKND2D0BWPHVT U610 ( .A1(N1330), .A2(N1293), .ZN(N123) );
  CKND2D0BWPHVT U611 ( .A1(N67), .A2(N1242), .ZN(N1227) );
  CKND2D0BWPHVT U612 ( .A1(N711), .A2(N130), .ZN(N1209) );
  CKND2D0BWPHVT U613 ( .A1(N1156), .A2(N383), .ZN(N130) );
  CKND2D0BWPHVT U614 ( .A1(N1605), .A2(N2), .ZN(N711) );
  CKND2D0BWPHVT U615 ( .A1(N203), .A2(N1813), .ZN(N1204) );
  CKND2D0BWPHVT U616 ( .A1(N605), .A2(N1091), .ZN(N1813) );
  CKND2D0BWPHVT U617 ( .A1(N462), .A2(N740), .ZN(N203) );
  ND3D0BWPHVT U618 ( .A1(n423), .A2(N326), .A3(N698), .ZN(N1190) );
  NR2D0BWPHVT U619 ( .A1(N1232), .A2(N229), .ZN(N698) );
  AN2D0BWPHVT U620 ( .A1(N142), .A2(N263), .Z(N1175) );
  CKND2D0BWPHVT U621 ( .A1(N864), .A2(N1556), .ZN(N263) );
  CKND2D0BWPHVT U622 ( .A1(N877), .A2(N1354), .ZN(N1556) );
  CKND0BWPHVT U623 ( .I(N1625), .ZN(N1354) );
  CKND2D0BWPHVT U624 ( .A1(N8), .A2(N1625), .ZN(N864) );
  CKND2D0BWPHVT U625 ( .A1(n419), .A2(N749), .ZN(N1625) );
  NR2D0BWPHVT U626 ( .A1(n424), .A2(N304), .ZN(n419) );
  CKND0BWPHVT U627 ( .I(N1283), .ZN(n424) );
  CKND2D0BWPHVT U628 ( .A1(N147), .A2(N390), .ZN(N1283) );
  CKND0BWPHVT U629 ( .I(N76), .ZN(N390) );
  CKND0BWPHVT U630 ( .I(N1087), .ZN(N147) );
  CKND2D0BWPHVT U631 ( .A1(N1502), .A2(N1077), .ZN(N142) );
  CKND2D0BWPHVT U632 ( .A1(N1577), .A2(N1074), .ZN(N1160) );
  ND3D0BWPHVT U633 ( .A1(N326), .A2(N1012), .A3(n423), .ZN(N1158) );
  AN3D0BWPHVT U634 ( .A1(N1429), .A2(N131), .A3(N1501), .Z(n423) );
  CKND0BWPHVT U635 ( .I(N1847), .ZN(N131) );
  CKND2D0BWPHVT U636 ( .A1(N402), .A2(N1332), .ZN(N1151) );
  CKND2D0BWPHVT U637 ( .A1(N1679), .A2(N389), .ZN(N1092) );
  CKND0BWPHVT U638 ( .I(N77), .ZN(N1077) );
  CKND2D0BWPHVT U639 ( .A1(N254), .A2(N925), .ZN(N1050) );
  CKND2D0BWPHVT U640 ( .A1(N943), .A2(N574), .ZN(N1033) );
  CKND2D0BWPHVT U641 ( .A1(N1130), .A2(N1021), .ZN(N574) );
  CKND2D0BWPHVT U642 ( .A1(N468), .A2(N1140), .ZN(N943) );
  CKND0BWPHVT U643 ( .I(N1130), .ZN(N1140) );
  CKND2D0BWPHVT U644 ( .A1(N1299), .A2(N1293), .ZN(N1130) );
  CKND2D0BWPHVT U645 ( .A1(N1087), .A2(N150), .ZN(N1025) );
  CKND2D0BWPHVT U646 ( .A1(n425), .A2(n426), .ZN(N1087) );
  NR4D0BWPHVT U647 ( .A1(N909), .A2(N462), .A3(N1230), .A4(N300), .ZN(n426) );
  CKND0BWPHVT U648 ( .I(N425), .ZN(N300) );
  ND3D0BWPHVT U649 ( .A1(N1146), .A2(N72), .A3(n427), .ZN(N425) );
  CKND0BWPHVT U650 ( .I(N605), .ZN(N462) );
  ND4D0BWPHVT U651 ( .A1(N1757), .A2(N341), .A3(n428), .A4(N630), .ZN(N605) );
  AN2D0BWPHVT U652 ( .A1(N1084), .A2(N264), .Z(n428) );
  CKND0BWPHVT U653 ( .I(N628), .ZN(N909) );
  ND3D0BWPHVT U654 ( .A1(N1641), .A2(N1501), .A3(n427), .ZN(N628) );
  NR4D0BWPHVT U655 ( .A1(N933), .A2(N1152), .A3(N1202), .A4(N728), .ZN(n425)
         );
  CKND0BWPHVT U656 ( .I(N1346), .ZN(N728) );
  ND3D0BWPHVT U657 ( .A1(N1641), .A2(N341), .A3(n429), .ZN(N1346) );
  CKND0BWPHVT U658 ( .I(N1477), .ZN(N1202) );
  ND3D0BWPHVT U659 ( .A1(N72), .A2(N1641), .A3(n429), .ZN(N1477) );
  CKND0BWPHVT U660 ( .I(N1587), .ZN(N1152) );
  ND3D0BWPHVT U661 ( .A1(N1146), .A2(N725), .A3(n429), .ZN(N1587) );
  AN3D0BWPHVT U662 ( .A1(N264), .A2(N1084), .A3(N1012), .Z(n429) );
  CKND0BWPHVT U663 ( .I(N402), .ZN(N933) );
  ND3D0BWPHVT U664 ( .A1(N1757), .A2(N341), .A3(n427), .ZN(N402) );
  CKND0BWPHVT U665 ( .I(N468), .ZN(N1021) );
  CKND2D0BWPHVT U666 ( .A1(N150), .A2(N76), .ZN(N468) );
  CKND2D0BWPHVT U667 ( .A1(n430), .A2(n431), .ZN(N76) );
  NR4D0BWPHVT U668 ( .A1(N727), .A2(N179), .A3(N743), .A4(N1156), .ZN(n431) );
  CKND0BWPHVT U669 ( .I(N1605), .ZN(N1156) );
  ND3D0BWPHVT U670 ( .A1(n432), .A2(N1429), .A3(N72), .ZN(N1605) );
  CKND0BWPHVT U671 ( .I(N1651), .ZN(N743) );
  ND3D0BWPHVT U672 ( .A1(N1501), .A2(n433), .A3(N1641), .ZN(N1651) );
  NR2D0BWPHVT U673 ( .A1(N1131), .A2(N762), .ZN(N1641) );
  CKND0BWPHVT U674 ( .I(N35), .ZN(N179) );
  ND3D0BWPHVT U675 ( .A1(n432), .A2(N1429), .A3(N341), .ZN(N35) );
  NR4D0BWPHVT U676 ( .A1(N712), .A2(N1679), .A3(N1763), .A4(N607), .ZN(n430)
         );
  CKND0BWPHVT U677 ( .I(N1161), .ZN(N1763) );
  ND3D0BWPHVT U678 ( .A1(N1501), .A2(n432), .A3(N1146), .ZN(N1161) );
  CKND0BWPHVT U679 ( .I(N117), .ZN(N1679) );
  ND3D0BWPHVT U680 ( .A1(N341), .A2(n433), .A3(N1146), .ZN(N117) );
  CKND0BWPHVT U681 ( .I(N1297), .ZN(N712) );
  ND3D0BWPHVT U682 ( .A1(N72), .A2(n433), .A3(N1146), .ZN(N1297) );
  NR2D0BWPHVT U683 ( .A1(N736), .A2(N1410), .ZN(N72) );
  CKND2D0BWPHVT U684 ( .A1(N564), .A2(N172), .ZN(N1006) );
  CKND2D0BWPHVT U685 ( .A1(N502), .A2(N1104), .ZN(N172) );
  CKND2D0BWPHVT U686 ( .A1(N727), .A2(N31), .ZN(N564) );
  CKND0BWPHVT U687 ( .I(N502), .ZN(N727) );
  ND3D0BWPHVT U688 ( .A1(N1429), .A2(n433), .A3(N725), .ZN(N502) );
  NR2D0BWPHVT U689 ( .A1(N1773), .A2(N736), .ZN(N725) );
  CKND0BWPHVT U690 ( .I(N414), .ZN(N736) );
  AN3D0BWPHVT U691 ( .A1(N264), .A2(N537), .A3(N630), .Z(n433) );
  NR2D0BWPHVT U692 ( .A1(N154), .A2(N1232), .ZN(N630) );
  NR2D0BWPHVT U693 ( .A1(N1113), .A2(N292), .ZN(N1429) );
  CKND2D0BWPHVT U694 ( .A1(N479), .A2(N1248), .ZN(N1004) );
  CKND2D0BWPHVT U695 ( .A1(N607), .A2(N1596), .ZN(N1248) );
  CKND0BWPHVT U696 ( .I(N1010), .ZN(N607) );
  CKND2D0BWPHVT U697 ( .A1(N1010), .A2(N1136), .ZN(N479) );
  ND3D0BWPHVT U698 ( .A1(N1501), .A2(n432), .A3(N1757), .ZN(N1010) );
  NR2D0BWPHVT U699 ( .A1(N762), .A2(N1113), .ZN(N1757) );
  CKND0BWPHVT U700 ( .I(N292), .ZN(N762) );
  AN3D0BWPHVT U701 ( .A1(N264), .A2(N537), .A3(N1012), .Z(n432) );
  CKND2D0BWPHVT U702 ( .A1(N1847), .A2(N1349), .ZN(N537) );
  ND3D0BWPHVT U703 ( .A1(n434), .A2(N1273), .A3(N1554), .ZN(N1349) );
  CKND0BWPHVT U704 ( .I(N1299), .ZN(n434) );
  CKND2D0BWPHVT U705 ( .A1(N1502), .A2(N1355), .ZN(N1299) );
  CKND0BWPHVT U706 ( .I(N1048), .ZN(N1355) );
  NR2D0BWPHVT U707 ( .A1(N1513), .A2(N1166), .ZN(N264) );
  CKND0BWPHVT U708 ( .I(N1063), .ZN(N1513) );
  NR2D0BWPHVT U709 ( .A1(N1410), .A2(N414), .ZN(N1501) );
  CKND2D0BWPHVT U710 ( .A1(N1230), .A2(N562), .ZN(N1000) );
  CKND0BWPHVT U711 ( .I(N59), .ZN(N1230) );
  ND3D0BWPHVT U712 ( .A1(N1146), .A2(N341), .A3(n427), .ZN(N59) );
  AN3D0BWPHVT U713 ( .A1(N1012), .A2(N1084), .A3(N326), .Z(n427) );
  NR2D0BWPHVT U714 ( .A1(N1166), .A2(N1063), .ZN(N326) );
  CKND2D0BWPHVT U715 ( .A1(N1826), .A2(N1447), .ZN(N1063) );
  CKND2D0BWPHVT U716 ( .A1(N1117), .A2(N344), .ZN(N1447) );
  CKND0BWPHVT U717 ( .I(N724), .ZN(N344) );
  CKND2D0BWPHVT U718 ( .A1(N724), .A2(N1282), .ZN(N1826) );
  CKND0BWPHVT U719 ( .I(N1117), .ZN(N1282) );
  CKND2D0BWPHVT U720 ( .A1(N226), .A2(N304), .ZN(N1117) );
  CKND2D0BWPHVT U721 ( .A1(N1692), .A2(N1038), .ZN(N226) );
  CKND2D0BWPHVT U722 ( .A1(N1330), .A2(N1300), .ZN(N1038) );
  CKND2D0BWPHVT U723 ( .A1(N938), .A2(N1293), .ZN(N1692) );
  CKND0BWPHVT U724 ( .I(N1300), .ZN(N1293) );
  CKND2D0BWPHVT U725 ( .A1(N487), .A2(N365), .ZN(N1300) );
  CKND2D0BWPHVT U726 ( .A1(N501), .A2(N93), .ZN(N365) );
  CKND0BWPHVT U727 ( .I(N24), .ZN(N93) );
  CKND0BWPHVT U728 ( .I(N1214), .ZN(N501) );
  CKND2D0BWPHVT U729 ( .A1(N24), .A2(N1214), .ZN(N487) );
  CKND2D0BWPHVT U730 ( .A1(N308), .A2(N244), .ZN(N1214) );
  CKND2D0BWPHVT U731 ( .A1(N1136), .A2(N31), .ZN(N244) );
  CKND2D0BWPHVT U732 ( .A1(N1104), .A2(N1596), .ZN(N308) );
  CKND2D0BWPHVT U733 ( .A1(N1838), .A2(N1823), .ZN(N24) );
  CKND2D0BWPHVT U734 ( .A1(N733), .A2(N423), .ZN(N1823) );
  CKND2D0BWPHVT U735 ( .A1(N751), .A2(N1406), .ZN(N1838) );
  CKND0BWPHVT U736 ( .I(N1330), .ZN(N938) );
  XNR2D0BWPHVT U737 ( .A1(N235), .A2(N1768), .ZN(N1330) );
  CKND2D0BWPHVT U738 ( .A1(N1053), .A2(N150), .ZN(N1768) );
  CKND0BWPHVT U739 ( .I(N1165), .ZN(N235) );
  CKND2D0BWPHVT U740 ( .A1(N685), .A2(N1561), .ZN(N1165) );
  CKND2D0BWPHVT U741 ( .A1(N841), .A2(N1091), .ZN(N1561) );
  CKND2D0BWPHVT U742 ( .A1(N1401), .A2(N740), .ZN(N685) );
  CKND2D0BWPHVT U743 ( .A1(N1126), .A2(N867), .ZN(N724) );
  CKND0BWPHVT U744 ( .I(N781), .ZN(N1166) );
  CKND2D0BWPHVT U745 ( .A1(N241), .A2(N867), .ZN(N781) );
  CKND2D0BWPHVT U746 ( .A1(N550), .A2(N304), .ZN(N867) );
  CKND2D0BWPHVT U747 ( .A1(N830), .A2(N1847), .ZN(N1084) );
  ND3D0BWPHVT U748 ( .A1(N77), .A2(N150), .A3(N1554), .ZN(N1847) );
  ND3D0BWPHVT U749 ( .A1(N1273), .A2(n435), .A3(N1554), .ZN(N830) );
  CKND2D0BWPHVT U750 ( .A1(N1134), .A2(N1653), .ZN(N1554) );
  CKND0BWPHVT U751 ( .I(N519), .ZN(n435) );
  CKND2D0BWPHVT U752 ( .A1(N1502), .A2(N1498), .ZN(N519) );
  CKND0BWPHVT U753 ( .I(N904), .ZN(N1498) );
  NR2D0BWPHVT U754 ( .A1(N191), .A2(N154), .ZN(N1012) );
  CKND0BWPHVT U755 ( .I(N229), .ZN(N154) );
  CKND2D0BWPHVT U756 ( .A1(N767), .A2(N961), .ZN(N229) );
  CKND0BWPHVT U757 ( .I(N1232), .ZN(N191) );
  CKND2D0BWPHVT U758 ( .A1(N1483), .A2(N1385), .ZN(N1232) );
  CKND2D0BWPHVT U759 ( .A1(N1118), .A2(N1812), .ZN(N1385) );
  CKND0BWPHVT U760 ( .I(N749), .ZN(N1812) );
  CKND2D0BWPHVT U761 ( .A1(N1549), .A2(N749), .ZN(N1483) );
  NR2D0BWPHVT U762 ( .A1(N1773), .A2(N414), .ZN(N341) );
  CKND2D0BWPHVT U763 ( .A1(N1544), .A2(N1452), .ZN(N414) );
  CKND2D0BWPHVT U764 ( .A1(N1511), .A2(N1869), .ZN(N1452) );
  CKND0BWPHVT U765 ( .I(N678), .ZN(N1869) );
  CKND0BWPHVT U766 ( .I(N1221), .ZN(N1511) );
  CKND2D0BWPHVT U767 ( .A1(N678), .A2(N1221), .ZN(N1544) );
  CKND2D0BWPHVT U768 ( .A1(N1408), .A2(N304), .ZN(N1221) );
  CKND2D0BWPHVT U769 ( .A1(N1163), .A2(N1090), .ZN(N1408) );
  CKND2D0BWPHVT U770 ( .A1(N611), .A2(N1016), .ZN(N1090) );
  CKND2D0BWPHVT U771 ( .A1(N11), .A2(N1189), .ZN(N1163) );
  CKND0BWPHVT U772 ( .I(N611), .ZN(N1189) );
  CKND2D0BWPHVT U773 ( .A1(N84), .A2(N375), .ZN(N611) );
  CKND2D0BWPHVT U774 ( .A1(N1154), .A2(N127), .ZN(N375) );
  CKND0BWPHVT U775 ( .I(N545), .ZN(N127) );
  CKND2D0BWPHVT U776 ( .A1(N545), .A2(N797), .ZN(N84) );
  CKND0BWPHVT U777 ( .I(N1154), .ZN(N797) );
  XNR2D0BWPHVT U778 ( .A1(N865), .A2(N1138), .ZN(N1154) );
  CKND0BWPHVT U779 ( .I(N486), .ZN(N865) );
  CKND2D0BWPHVT U780 ( .A1(N366), .A2(N1584), .ZN(N486) );
  CKND2D0BWPHVT U781 ( .A1(N416), .A2(N534), .ZN(N1584) );
  CKND2D0BWPHVT U782 ( .A1(N1670), .A2(N67), .ZN(N366) );
  XNR2D0BWPHVT U783 ( .A1(N310), .A2(N383), .ZN(N545) );
  CKND0BWPHVT U784 ( .I(N810), .ZN(N310) );
  CKND2D0BWPHVT U785 ( .A1(N1770), .A2(N1322), .ZN(N810) );
  CKND2D0BWPHVT U786 ( .A1(N513), .A2(N31), .ZN(N1322) );
  CKND2D0BWPHVT U787 ( .A1(N1104), .A2(N520), .ZN(N1770) );
  CKND0BWPHVT U788 ( .I(N1016), .ZN(N11) );
  ND3D0BWPHVT U789 ( .A1(N1134), .A2(N150), .A3(N328), .ZN(N1016) );
  CKND0BWPHVT U790 ( .I(N1410), .ZN(N1773) );
  CKND2D0BWPHVT U791 ( .A1(N873), .A2(N79), .ZN(N1410) );
  CKND2D0BWPHVT U792 ( .A1(N949), .A2(N510), .ZN(N79) );
  CKND2D0BWPHVT U793 ( .A1(N1142), .A2(N166), .ZN(N873) );
  CKND0BWPHVT U794 ( .I(N949), .ZN(N166) );
  CKND0BWPHVT U795 ( .I(N510), .ZN(N1142) );
  CKND2D0BWPHVT U796 ( .A1(N234), .A2(N304), .ZN(N510) );
  CKND2D0BWPHVT U797 ( .A1(N56), .A2(N1661), .ZN(N234) );
  CKND2D0BWPHVT U798 ( .A1(N1315), .A2(N378), .ZN(N1661) );
  CKND2D0BWPHVT U799 ( .A1(N1257), .A2(N367), .ZN(N56) );
  CKND0BWPHVT U800 ( .I(N378), .ZN(N367) );
  XNR2D0BWPHVT U801 ( .A1(N783), .A2(N1331), .ZN(N378) );
  CKND0BWPHVT U802 ( .I(N1800), .ZN(N783) );
  CKND2D0BWPHVT U803 ( .A1(N49), .A2(N232), .ZN(N1800) );
  CKND2D0BWPHVT U804 ( .A1(N124), .A2(N31), .ZN(N232) );
  CKND0BWPHVT U805 ( .I(N1104), .ZN(N31) );
  CKND2D0BWPHVT U806 ( .A1(N1104), .A2(N389), .ZN(N49) );
  CKND0BWPHVT U807 ( .I(N1315), .ZN(N1257) );
  XNR2D0BWPHVT U808 ( .A1(N1237), .A2(N1479), .ZN(N1315) );
  CKND0BWPHVT U809 ( .I(N568), .ZN(N1237) );
  CKND2D0BWPHVT U810 ( .A1(N1133), .A2(N1065), .ZN(N568) );
  CKND2D0BWPHVT U811 ( .A1(N412), .A2(N227), .ZN(N1065) );
  CKND0BWPHVT U812 ( .I(N518), .ZN(N412) );
  CKND2D0BWPHVT U813 ( .A1(N518), .A2(N562), .ZN(N1133) );
  XNR2D0BWPHVT U814 ( .A1(N206), .A2(N67), .ZN(N518) );
  CKND0BWPHVT U815 ( .I(N1242), .ZN(N206) );
  ND3D0BWPHVT U816 ( .A1(N150), .A2(N550), .A3(N241), .ZN(N1242) );
  NR2D0BWPHVT U817 ( .A1(N1131), .A2(N292), .ZN(N1146) );
  CKND2D0BWPHVT U818 ( .A1(N922), .A2(N242), .ZN(N292) );
  CKND2D0BWPHVT U819 ( .A1(N1320), .A2(N935), .ZN(N242) );
  CKND0BWPHVT U820 ( .I(N330), .ZN(N935) );
  CKND2D0BWPHVT U821 ( .A1(N330), .A2(N174), .ZN(N922) );
  CKND0BWPHVT U822 ( .I(N1320), .ZN(N174) );
  CKND2D0BWPHVT U823 ( .A1(N328), .A2(N961), .ZN(N1320) );
  CKND2D0BWPHVT U824 ( .A1(N1134), .A2(N304), .ZN(N961) );
  CKND2D0BWPHVT U825 ( .A1(N304), .A2(N1179), .ZN(N330) );
  CKND2D0BWPHVT U826 ( .A1(N88), .A2(N152), .ZN(N1179) );
  CKND2D0BWPHVT U827 ( .A1(N1819), .A2(N1672), .ZN(N152) );
  CKND0BWPHVT U828 ( .I(N1748), .ZN(N1672) );
  CKND2D0BWPHVT U829 ( .A1(N823), .A2(N1748), .ZN(N88) );
  CKND2D0BWPHVT U830 ( .A1(N548), .A2(N276), .ZN(N1748) );
  CKND2D0BWPHVT U831 ( .A1(N1756), .A2(N1479), .ZN(N276) );
  CKND0BWPHVT U832 ( .I(N884), .ZN(N1479) );
  CKND2D0BWPHVT U833 ( .A1(N884), .A2(N64), .ZN(N548) );
  CKND0BWPHVT U834 ( .I(N1756), .ZN(N64) );
  XNR2D0BWPHVT U835 ( .A1(N1015), .A2(N1596), .ZN(N1756) );
  CKND0BWPHVT U836 ( .I(N870), .ZN(N1015) );
  CKND2D0BWPHVT U837 ( .A1(N1717), .A2(N1172), .ZN(N870) );
  CKND2D0BWPHVT U838 ( .A1(N1670), .A2(N979), .ZN(N1172) );
  CKND2D0BWPHVT U839 ( .A1(N1405), .A2(N534), .ZN(N1717) );
  XNR2D0BWPHVT U840 ( .A1(N684), .A2(N288), .ZN(N884) );
  CKND2D0BWPHVT U841 ( .A1(N223), .A2(N1602), .ZN(N288) );
  CKND2D0BWPHVT U842 ( .A1(N1091), .A2(N800), .ZN(N1602) );
  CKND2D0BWPHVT U843 ( .A1(N1332), .A2(N740), .ZN(N223) );
  CKND0BWPHVT U844 ( .I(N1091), .ZN(N740) );
  CKND0BWPHVT U845 ( .I(N1819), .ZN(N823) );
  XNR2D0BWPHVT U846 ( .A1(N1577), .A2(N984), .ZN(N1819) );
  CKND0BWPHVT U847 ( .I(N626), .ZN(N1577) );
  ND3D0BWPHVT U848 ( .A1(N1134), .A2(N150), .A3(N767), .ZN(N626) );
  CKND0BWPHVT U849 ( .I(N1113), .ZN(N1131) );
  CKND2D0BWPHVT U850 ( .A1(N1600), .A2(N1099), .ZN(N1113) );
  CKND2D0BWPHVT U851 ( .A1(N1115), .A2(N1522), .ZN(N1099) );
  CKND0BWPHVT U852 ( .I(N882), .ZN(N1522) );
  CKND0BWPHVT U853 ( .I(N1047), .ZN(N1115) );
  CKND2D0BWPHVT U854 ( .A1(N1047), .A2(N882), .ZN(N1600) );
  CKND2D0BWPHVT U855 ( .A1(N304), .A2(N29), .ZN(N1047) );
  CKND2D0BWPHVT U856 ( .A1(N757), .A2(N1699), .ZN(N29) );
  CKND2D0BWPHVT U857 ( .A1(N1362), .A2(N544), .ZN(N1699) );
  CKND0BWPHVT U858 ( .I(N824), .ZN(N544) );
  CKND0BWPHVT U859 ( .I(N258), .ZN(N1362) );
  CKND2D0BWPHVT U860 ( .A1(N258), .A2(N824), .ZN(N757) );
  CKND2D0BWPHVT U861 ( .A1(N707), .A2(N408), .ZN(N824) );
  CKND2D0BWPHVT U862 ( .A1(N1406), .A2(N744), .ZN(N408) );
  CKND2D0BWPHVT U863 ( .A1(N733), .A2(N1664), .ZN(N707) );
  CKND0BWPHVT U864 ( .I(N744), .ZN(N1664) );
  CKND2D0BWPHVT U865 ( .A1(N955), .A2(N1309), .ZN(N744) );
  CKND2D0BWPHVT U866 ( .A1(N1401), .A2(N1711), .ZN(N1309) );
  CKND2D0BWPHVT U867 ( .A1(N841), .A2(N1359), .ZN(N955) );
  CKND0BWPHVT U868 ( .I(N1406), .ZN(N733) );
  XNR2D0BWPHVT U869 ( .A1(N954), .A2(N389), .ZN(N1406) );
  CKND0BWPHVT U870 ( .I(N124), .ZN(N389) );
  CKND0BWPHVT U871 ( .I(N1667), .ZN(N954) );
  CKND2D0BWPHVT U872 ( .A1(N623), .A2(N1685), .ZN(N1667) );
  CKND2D0BWPHVT U873 ( .A1(N513), .A2(N979), .ZN(N1685) );
  CKND0BWPHVT U874 ( .I(N1405), .ZN(N979) );
  CKND2D0BWPHVT U875 ( .A1(N1405), .A2(N520), .ZN(N623) );
  CKND0BWPHVT U876 ( .I(N513), .ZN(N520) );
  XNR2D0BWPHVT U877 ( .A1(N1011), .A2(N254), .ZN(N258) );
  CKND0BWPHVT U878 ( .I(N925), .ZN(N1011) );
  ND3D0BWPHVT U879 ( .A1(N150), .A2(N550), .A3(N1126), .ZN(N925) );
  CKND0BWPHVT U880 ( .I(N1653), .ZN(N550) );
  CKND0BWPHVT U881 ( .I(N1549), .ZN(N1118) );
  CKND2D0BWPHVT U882 ( .A1(N8), .A2(N304), .ZN(N1549) );
  CKND0BWPHVT U883 ( .I(N1273), .ZN(N304) );
  CKND0BWPHVT U884 ( .I(N877), .ZN(N8) );
  XNR2D0BWPHVT U885 ( .A1(N911), .A2(N1507), .ZN(N877) );
  CKND2D0BWPHVT U886 ( .A1(N972), .A2(N415), .ZN(N1507) );
  CKND2D0BWPHVT U887 ( .A1(N939), .A2(N1687), .ZN(N415) );
  CKND2D0BWPHVT U888 ( .A1(N1066), .A2(N63), .ZN(N972) );
  CKND0BWPHVT U889 ( .I(N939), .ZN(N63) );
  CKND2D0BWPHVT U890 ( .A1(N1239), .A2(N1218), .ZN(N939) );
  CKND2D0BWPHVT U891 ( .A1(N1136), .A2(N800), .ZN(N1218) );
  CKND0BWPHVT U892 ( .I(N1332), .ZN(N800) );
  CKND2D0BWPHVT U893 ( .A1(N1332), .A2(N1596), .ZN(N1239) );
  CKND0BWPHVT U894 ( .I(N1136), .ZN(N1596) );
  CKND0BWPHVT U895 ( .I(N1687), .ZN(N1066) );
  CKND2D0BWPHVT U896 ( .A1(N1141), .A2(N150), .ZN(N1687) );
  CKND0BWPHVT U897 ( .I(N1502), .ZN(N150) );
  CKND0BWPHVT U898 ( .I(N1767), .ZN(N911) );
  CKND2D0BWPHVT U899 ( .A1(N1491), .A2(N1127), .ZN(N1767) );
  CKND2D0BWPHVT U900 ( .A1(N673), .A2(N1359), .ZN(N1127) );
  CKND2D0BWPHVT U901 ( .A1(N1711), .A2(N1246), .ZN(N1491) );
  CKND0BWPHVT U902 ( .I(N673), .ZN(N1246) );
  CKND2D0BWPHVT U903 ( .A1(N52), .A2(N1277), .ZN(N673) );
  CKND2D0BWPHVT U904 ( .A1(N751), .A2(N841), .ZN(N1277) );
  CKND2D0BWPHVT U905 ( .A1(N423), .A2(N1401), .ZN(N52) );
  CKND0BWPHVT U906 ( .I(N841), .ZN(N1401) );
  XNR2D0BWPHVT U907 ( .A1(N660), .A2(N534), .ZN(N841) );
  CKND0BWPHVT U908 ( .I(N1670), .ZN(N534) );
  CKND0BWPHVT U909 ( .I(N1722), .ZN(N660) );
  CKND2D0BWPHVT U910 ( .A1(N42), .A2(N1662), .ZN(N1722) );
  CKND2D0BWPHVT U911 ( .A1(N416), .A2(N811), .ZN(N1662) );
  CKND0BWPHVT U912 ( .I(N684), .ZN(N811) );
  CKND2D0BWPHVT U913 ( .A1(N684), .A2(N67), .ZN(N42) );
  CKND0BWPHVT U914 ( .I(N416), .ZN(N67) );
  CKND0BWPHVT U915 ( .I(N751), .ZN(N423) );
  XNR2D0BWPHVT U916 ( .A1(N1123), .A2(N254), .ZN(N751) );
  CKND0BWPHVT U917 ( .I(N249), .ZN(N254) );
  CKND0BWPHVT U918 ( .I(N621), .ZN(N1123) );
  CKND2D0BWPHVT U919 ( .A1(N1714), .A2(N102), .ZN(N621) );
  CKND2D0BWPHVT U920 ( .A1(N287), .A2(N383), .ZN(N102) );
  CKND0BWPHVT U921 ( .I(N2), .ZN(N383) );
  CKND2D0BWPHVT U922 ( .A1(N2), .A2(N1331), .ZN(N1714) );
  CKND0BWPHVT U923 ( .I(N287), .ZN(N1331) );
  CKND0BWPHVT U924 ( .I(N1359), .ZN(N1711) );
  CKND2D0BWPHVT U925 ( .A1(N74), .A2(N732), .ZN(N1359) );
  CKND2D0BWPHVT U926 ( .A1(N1159), .A2(N227), .ZN(N732) );
  CKND2D0BWPHVT U927 ( .A1(N1766), .A2(N562), .ZN(N74) );
  CKND0BWPHVT U928 ( .I(N227), .ZN(N562) );
  CKND0BWPHVT U929 ( .I(N1159), .ZN(N1766) );
  CKND2D0BWPHVT U930 ( .A1(N1648), .A2(N1205), .ZN(N1159) );
  CKND2D0BWPHVT U931 ( .A1(N528), .A2(N984), .ZN(N1205) );
  CKND0BWPHVT U932 ( .I(N1074), .ZN(N984) );
  CKND2D0BWPHVT U933 ( .A1(N1074), .A2(N1138), .ZN(N1648) );
  CKND0BWPHVT U934 ( .I(N528), .ZN(N1138) );
endmodule

