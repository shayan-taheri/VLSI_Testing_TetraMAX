
module HFC2 (N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670, N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873);

input N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670;
output N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873;
  wire   N1622, N716, N1872, N873, N933, N1316, N1674, N1416, N1249, N305,
         N1698, N2, N77, N124, N227, N249, N287, N416, N513, N528, N678, N684,
         N749, N882, N949, N1074, N1091, N1104, N1134, N1136, N1273, N1332,
         N1405, N1502, N1670, N1042, N1722, N121, N785, N1241, N1383, N1569,
         N64, N1454, N386, N292, N1399, N315, N157, N1169, N229, N903, N389,
         N13, N569, N743, N270, N899, N681, N1257, N1407, N224, N1287, N676,
         N456, N1052, N813, N78, N364, N149, N7, N530, N1777, N1688, N981,
         N948, N266, N1609, N1326, N1536, N1501, N967, N50, N567, N538, N481,
         N1029, N212, N883, N698, N602, N163, N1404, N831, N288, N1763, N952,
         N437, N745, N334, N1166, N21, N1366, N777, N462, N95, N649, N648,
         N144, N24, N319, N609, N1096, N932, N909, N449, N181, N1408, N438,
         N566, N790, N652, N761, N401, N906, N52, N852, N519, N726, N258,
         N1751, N441, N263, N531, N268, N1197, N276, N654, N1759, N911, N543,
         N1479, N1195, N580, N1388, N1030, N1253, N90, N1248, N1786, N837,
         N1431, N1039, N550, N1799, N1244, N997, N1470, N668, N1682, N717,
         N1518, N1014, N941, N1508, N593, N637, N500, N582, N751, N1238, N1562,
         N1100, N1499, N812, N271, N409, N910, N669, N1789, N1769, N486, N1748,
         N1398, N1276, N562, N1066, N402, N505, N1060, N1665, N841, N973, N92,
         N1409, N591, N1511, N650, N969, N109, N1440, N1775, N1112, N205, N256,
         N670, N1321, N1595, N311, N1328, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440;
  assign N1346 = N1622;
  assign N700 = N716;
  assign N920 = N1872;
  assign N417 = N873;
  assign N559 = N933;
  assign N1133 = N1316;
  assign N342 = N1674;
  assign N439 = N1416;
  assign N539 = N1249;
  assign N1863 = N305;
  assign N1746 = N305;
  assign N380 = N305;
  assign N91 = N305;
  assign N247 = N1698;
  assign N617 = N1698;
  assign N130 = N1698;
  assign N284 = N1698;
  assign N350 = N1698;
  assign N1119 = N1698;
  assign N1761 = N2;
  assign N619 = N2;
  assign N388 = N2;
  assign N278 = N2;
  assign N1385 = N77;
  assign N1258 = N124;
  assign N1842 = N124;
  assign N521 = N124;
  assign N203 = N124;
  assign N620 = N227;
  assign N1788 = N227;
  assign N1114 = N227;
  assign N1079 = N227;
  assign N1334 = N249;
  assign N1159 = N249;
  assign N988 = N249;
  assign N455 = N249;
  assign N367 = N249;
  assign N423 = N287;
  assign N1468 = N287;
  assign N878 = N287;
  assign N335 = N287;
  assign N281 = N416;
  assign N1638 = N416;
  assign N1584 = N416;
  assign N1504 = N416;
  assign N190 = N416;
  assign N67 = N513;
  assign N171 = N513;
  assign N20 = N513;
  assign N11 = N513;
  assign N553 = N528;
  assign N369 = N528;
  assign N156 = N528;
  assign N81 = N528;
  assign N1430 = N678;
  assign N817 = N678;
  assign N1568 = N684;
  assign N1672 = N684;
  assign N1546 = N684;
  assign N816 = N684;
  assign N166 = N684;
  assign N1345 = N749;
  assign N17 = N749;
  assign N666 = N882;
  assign N546 = N882;
  assign N1652 = N949;
  assign N452 = N949;
  assign N810 = N1074;
  assign N1826 = N1074;
  assign N712 = N1074;
  assign N696 = N1074;
  assign N937 = N1091;
  assign N1767 = N1091;
  assign N800 = N1091;
  assign N799 = N1091;
  assign N770 = N1091;
  assign N482 = N1091;
  assign N1530 = N1104;
  assign N1510 = N1104;
  assign N604 = N1104;
  assign N45 = N1104;
  assign N795 = N1134;
  assign N738 = N1134;
  assign N1681 = N1136;
  assign N1008 = N1136;
  assign N847 = N1136;
  assign N460 = N1136;
  assign N225 = N1136;
  assign N1118 = N1273;
  assign N688 = N1273;
  assign N1363 = N1332;
  assign N1450 = N1332;
  assign N970 = N1332;
  assign N956 = N1332;
  assign N551 = N1332;
  assign N80 = N1332;
  assign N1433 = N1405;
  assign N850 = N1405;
  assign N636 = N1405;
  assign N143 = N1405;
  assign N1785 = N1502;
  assign N1588 = N1502;
  assign N1532 = N1502;
  assign N820 = N1670;
  assign N1534 = N1670;
  assign N1339 = N1670;
  assign N375 = N1670;
  assign N96 = N1670;
  assign N1675 = N1042;
  assign N834 = N1042;
  assign N1379 = N1722;
  assign N931 = N1722;
  assign N1571 = N121;
  assign N748 = N121;
  assign N239 = N121;
  assign N374 = N121;
  assign N356 = N785;
  assign N301 = N785;
  assign N639 = N1241;
  assign N951 = N1383;
  assign N410 = N1569;
  assign N1041 = N1569;
  assign N775 = N64;
  assign N1349 = N1454;
  assign N74 = N1454;
  assign N1246 = N1454;
  assign N869 = N1454;
  assign N405 = N1454;
  assign N856 = N386;
  assign N1325 = N292;
  assign N420 = N292;
  assign N1648 = N1399;
  assign N890 = N315;
  assign N297 = N157;
  assign N384 = N1169;
  assign N1774 = N229;
  assign N783 = N229;
  assign N1097 = N903;
  assign N1056 = N389;
  assign N1716 = N13;
  assign N1654 = N13;
  assign N805 = N13;
  assign N261 = N13;
  assign N231 = N13;
  assign N444 = N569;
  assign N1493 = N743;
  assign N979 = N270;
  assign N308 = N270;
  assign N1464 = N899;
  assign N1111 = N899;
  assign N905 = N899;
  assign N809 = N899;
  assign N1642 = N681;
  assign N1009 = N681;
  assign N893 = N681;
  assign N661 = N681;
  assign N1377 = N681;
  assign N1080 = N1257;
  assign N1639 = N1407;
  assign N975 = N1407;
  assign N1712 = N224;
  assign N1151 = N1287;
  assign N989 = N1287;
  assign N140 = N1287;
  assign N324 = N1287;
  assign N830 = N1287;
  assign N1723 = N676;
  assign N446 = N676;
  assign N1825 = N456;
  assign N1188 = N456;
  assign N996 = N456;
  assign N927 = N456;
  assign N889 = N456;
  assign N468 = N1052;
  assign N1662 = N813;
  assign N244 = N813;
  assign N104 = N813;
  assign N58 = N813;
  assign N48 = N813;
  assign N1286 = N813;
  assign N1815 = N78;
  assign N1796 = N78;
  assign N1362 = N78;
  assign N443 = N78;
  assign N914 = N78;
  assign N1664 = N364;
  assign N947 = N149;
  assign N394 = N149;
  assign N1634 = N7;
  assign N491 = N7;
  assign N732 = N530;
  assign N1780 = N1777;
  assign N597 = N1777;
  assign N245 = N1777;
  assign N213 = N1777;
  assign N861 = N1777;
  assign N218 = N1777;
  assign N1089 = N1777;
  assign N360 = N1777;
  assign N1602 = N1688;
  assign N1218 = N981;
  assign N1182 = N981;
  assign N435 = N981;
  assign N155 = N981;
  assign N122 = N981;
  assign N798 = N981;
  assign N1491 = N948;
  assign N1607 = N266;
  assign N1498 = N266;
  assign N1063 = N266;
  assign N433 = N266;
  assign N131 = N266;
  assign N1463 = N1609;
  assign N1819 = N1326;
  assign N1485 = N1326;
  assign N1304 = N1326;
  assign N16 = N1326;
  assign N1717 = N1326;
  assign N1201 = N1536;
  assign N250 = N1536;
  assign N1572 = N1501;
  assign N1553 = N1501;
  assign N912 = N1501;
  assign N832 = N1501;
  assign N264 = N1501;
  assign N1772 = N1501;
  assign N757 = N967;
  assign N1870 = N50;
  assign N1747 = N50;
  assign N1342 = N567;
  assign N1291 = N538;
  assign N66 = N538;
  assign N223 = N481;
  assign N1168 = N1029;
  assign N731 = N1029;
  assign N1022 = N212;
  assign N958 = N212;
  assign N699 = N883;
  assign N611 = N883;
  assign N1856 = N698;
  assign N1288 = N698;
  assign N98 = N698;
  assign N1012 = N698;
  assign N1 = N602;
  assign N671 = N602;
  assign N1694 = N163;
  assign N844 = N163;
  assign N771 = N163;
  assign N759 = N163;
  assign N291 = N163;
  assign N129 = N163;
  assign N1770 = N163;
  assign N1301 = N1404;
  assign N1262 = N1404;
  assign N483 = N831;
  assign N285 = N831;
  assign N93 = N831;
  assign N1154 = N831;
  assign N373 = N288;
  assign N202 = N288;
  assign N875 = N1763;
  assign N1261 = N1763;
  assign N1092 = N952;
  assign N83 = N437;
  assign N1378 = N745;
  assign N1170 = N745;
  assign N1123 = N745;
  assign N913 = N745;
  assign N925 = N745;
  assign N859 = N334;
  assign N1153 = N1166;
  assign N746 = N1166;
  assign N404 = N21;
  assign N788 = N1366;
  assign N641 = N1366;
  assign N479 = N1366;
  assign N338 = N1366;
  assign N312 = N1366;
  assign N272 = N1366;
  assign N238 = N1366;
  assign N1587 = N1366;
  assign N1800 = N777;
  assign N1226 = N777;
  assign N1161 = N777;
  assign N1392 = N777;
  assign N1585 = N462;
  assign N1269 = N462;
  assign N522 = N462;
  assign N1163 = N95;
  assign N1200 = N649;
  assign N826 = N649;
  assign N414 = N649;
  assign N359 = N649;
  assign N6 = N649;
  assign N153 = N649;
  assign N1350 = N648;
  assign N1419 = N144;
  assign N667 = N24;
  assign N833 = N319;
  assign N984 = N609;
  assign N383 = N1096;
  assign N578 = N932;
  assign N495 = N909;
  assign N1138 = N449;
  assign N1846 = N181;
  assign N325 = N1408;
  assign N1084 = N438;
  assign N1471 = N566;
  assign N59 = N790;
  assign N86 = N652;
  assign N1023 = N761;
  assign N188 = N761;
  assign N585 = N401;
  assign N1847 = N906;
  assign N675 = N52;
  assign N968 = N852;
  assign N1415 = N519;
  assign N279 = N726;
  assign N277 = N726;
  assign N1297 = N258;
  assign N588 = N1751;
  assign N1848 = N441;
  assign N317 = N263;
  assign N170 = N531;
  assign N576 = N268;
  assign N178 = N1197;
  assign N217 = N276;
  assign N1538 = N654;
  assign N1641 = N1759;
  assign N430 = N911;
  assign N1446 = N543;
  assign N1315 = N1479;
  assign N79 = N1195;
  assign N603 = N580;
  assign N1497 = N580;
  assign N262 = N580;
  assign N1237 = N1388;
  assign N1494 = N1030;
  assign N100 = N1253;
  assign N827 = N90;
  assign N990 = N1248;
  assign N322 = N1786;
  assign N145 = N837;
  assign N1002 = N1431;
  assign N864 = N1431;
  assign N1110 = N1431;
  assign N151 = N1431;
  assign N209 = N1431;
  assign N564 = N1039;
  assign N640 = N550;
  assign N605 = N1799;
  assign N211 = N1799;
  assign N25 = N1244;
  assign N557 = N997;
  assign N1324 = N1470;
  assign N1072 = N1470;
  assign N982 = N668;
  assign N139 = N1682;
  assign N1338 = N1682;
  assign N631 = N717;
  assign N160 = N1518;
  assign N112 = N1014;
  assign N1857 = N941;
  assign N1624 = N941;
  assign N1216 = N1508;
  assign N545 = N1508;
  assign N1320 = N593;
  assign N330 = N593;
  assign N1728 = N637;
  assign N1678 = N500;
  assign N436 = N582;
  assign N1484 = N751;
  assign N1813 = N751;
  assign N892 = N1238;
  assign N536 = N1562;
  assign N280 = N1100;
  assign N422 = N1100;
  assign N714 = N1499;
  assign N103 = N812;
  assign N1278 = N271;
  assign N126 = N271;
  assign N29 = N409;
  assign N626 = N910;
  assign N629 = N669;
  assign N1547 = N1789;
  assign N1214 = N1769;
  assign N345 = N1769;
  assign N318 = N1769;
  assign N1145 = N1769;
  assign N1749 = N1769;
  assign N204 = N1769;
  assign N294 = N1769;
  assign N403 = N1769;
  assign N526 = N1769;
  assign N307 = N486;
  assign N61 = N1748;
  assign N1418 = N1398;
  assign N821 = N1276;
  assign N1228 = N562;
  assign N198 = N1066;
  assign N363 = N402;
  assign N469 = N505;
  assign N31 = N1060;
  assign N1563 = N1665;
  assign N1567 = N841;
  assign N1083 = N973;
  assign N894 = N973;
  assign N794 = N92;
  assign N1805 = N1409;
  assign N901 = N591;
  assign N186 = N1511;
  assign N33 = N650;
  assign N1421 = N650;
  assign N159 = N650;
  assign N908 = N969;
  assign N735 = N969;
  assign N1353 = N109;
  assign N517 = N109;
  assign N634 = N1440;
  assign N219 = N1440;
  assign N560 = N1775;
  assign N1684 = N1775;
  assign N659 = N1112;
  assign N87 = N205;
  assign N41 = N205;
  assign N838 = N256;
  assign N174 = N670;
  assign N1808 = N1321;
  assign N117 = N1595;
  assign N709 = N311;
  assign N1047 = N1328;

  AN2D0BWPHVT U477 ( .A1(N13), .A2(N615), .Z(N97) );
  CKND2D0BWPHVT U478 ( .A1(N1249), .A2(N883), .ZN(N910) );
  NR2D0BWPHVT U479 ( .A1(N1156), .A2(N1088), .ZN(N891) );
  CKND0BWPHVT U480 ( .I(N1511), .ZN(N883) );
  CKND2D0BWPHVT U481 ( .A1(N1416), .A2(N1447), .ZN(N881) );
  CKND2D0BWPHVT U482 ( .A1(N952), .A2(N315), .ZN(N852) );
  CKND0BWPHVT U483 ( .I(N205), .ZN(N952) );
  CKND2D0BWPHVT U484 ( .A1(N267), .A2(N1443), .ZN(N824) );
  CKND2D0BWPHVT U485 ( .A1(N1478), .A2(N2), .ZN(N815) );
  CKND2D0BWPHVT U486 ( .A1(N981), .A2(N1210), .ZN(N808) );
  CKND2D0BWPHVT U487 ( .A1(N862), .A2(N973), .ZN(N807) );
  CKND2D0BWPHVT U488 ( .A1(N1371), .A2(N1327), .ZN(N787) );
  CKND2D0BWPHVT U489 ( .A1(N72), .A2(N1627), .ZN(N740) );
  CKND2D0BWPHVT U490 ( .A1(N1667), .A2(N649), .ZN(N72) );
  CKND2D0BWPHVT U491 ( .A1(N676), .A2(N602), .ZN(N674) );
  CKND2D0BWPHVT U492 ( .A1(N1769), .A2(N1091), .ZN(N669) );
  CKND2D0BWPHVT U493 ( .A1(N899), .A2(N676), .ZN(N668) );
  CKND2D0BWPHVT U494 ( .A1(N286), .A2(N236), .ZN(N664) );
  CKND2D0BWPHVT U495 ( .A1(N1169), .A2(N813), .ZN(N654) );
  CKND2D0BWPHVT U496 ( .A1(N1060), .A2(N227), .ZN(N637) );
  CKND2D0BWPHVT U497 ( .A1(N682), .A2(N1137), .ZN(N615) );
  CKND2D0BWPHVT U498 ( .A1(N1373), .A2(N751), .ZN(N682) );
  CKND0BWPHVT U499 ( .I(N530), .ZN(N1249) );
  CKND2D0BWPHVT U500 ( .A1(N941), .A2(N1431), .ZN(N550) );
  CKND2D0BWPHVT U501 ( .A1(N358), .A2(N481), .ZN(N549) );
  CKND2D0BWPHVT U502 ( .A1(N698), .A2(N15), .ZN(N542) );
  CKND2D0BWPHVT U503 ( .A1(N726), .A2(N205), .ZN(N519) );
  AN2D0BWPHVT U504 ( .A1(N13), .A2(N116), .Z(N510) );
  CKND2D0BWPHVT U505 ( .A1(N1609), .A2(N456), .ZN(N500) );
  CKND2D0BWPHVT U506 ( .A1(N82), .A2(N638), .ZN(N466) );
  CKND2D0BWPHVT U507 ( .A1(N1316), .A2(N1569), .ZN(N464) );
  CKND2D0BWPHVT U508 ( .A1(N234), .A2(N137), .ZN(N431) );
  CKND2D0BWPHVT U509 ( .A1(N393), .A2(N1606), .ZN(N413) );
  CKND2D0BWPHVT U510 ( .A1(N530), .A2(N1511), .ZN(N409) );
  CKND2D0BWPHVT U511 ( .A1(N302), .A2(N1355), .ZN(N393) );
  AN2D0BWPHVT U512 ( .A1(N13), .A2(N195), .Z(N387) );
  CKND2D0BWPHVT U513 ( .A1(N707), .A2(N1344), .ZN(N378) );
  CKND2D0BWPHVT U514 ( .A1(N323), .A2(N1326), .ZN(N707) );
  CKND2D0BWPHVT U515 ( .A1(N1095), .A2(N416), .ZN(N371) );
  CKND2D0BWPHVT U516 ( .A1(N1113), .A2(N496), .ZN(N362) );
  CKND2D0BWPHVT U517 ( .A1(N1142), .A2(N745), .ZN(N36) );
  CKND0BWPHVT U518 ( .I(N82), .ZN(N358) );
  CKND2D0BWPHVT U519 ( .A1(N1003), .A2(N121), .ZN(N357) );
  CKND2D0BWPHVT U520 ( .A1(N686), .A2(N570), .ZN(N34) );
  CKND2D0BWPHVT U521 ( .A1(N566), .A2(N249), .ZN(N570) );
  CKND2D0BWPHVT U522 ( .A1(N26), .A2(N813), .ZN(N686) );
  CKND2D0BWPHVT U523 ( .A1(N1742), .A2(N1458), .ZN(N300) );
  CKND2D0BWPHVT U524 ( .A1(N1683), .A2(N78), .ZN(N286) );
  CKND2D0BWPHVT U525 ( .A1(N633), .A2(N121), .ZN(N267) );
  CKND2D0BWPHVT U526 ( .A1(N181), .A2(N287), .ZN(N236) );
  CKND2D0BWPHVT U527 ( .A1(N660), .A2(N777), .ZN(N234) );
  CKND2D0BWPHVT U528 ( .A1(N450), .A2(N347), .ZN(N195) );
  CKND2D0BWPHVT U529 ( .A1(N52), .A2(N370), .ZN(N347) );
  CKND2D0BWPHVT U530 ( .A1(N502), .A2(N1512), .ZN(N450) );
  CKND0BWPHVT U531 ( .I(N370), .ZN(N502) );
  CKND2D0BWPHVT U532 ( .A1(n424), .A2(N678), .ZN(N370) );
  CKND2D0BWPHVT U533 ( .A1(N650), .A2(N941), .ZN(N1837) );
  CKND2D0BWPHVT U534 ( .A1(N1777), .A2(N163), .ZN(N1789) );
  CKND2D0BWPHVT U535 ( .A1(N911), .A2(N249), .ZN(N1759) );
  CKND2D0BWPHVT U536 ( .A1(N1460), .A2(N416), .ZN(N1742) );
  CKND0BWPHVT U537 ( .I(N941), .ZN(N676) );
  CKND2D0BWPHVT U538 ( .A1(N193), .A2(N528), .ZN(N1704) );
  CKND2D0BWPHVT U539 ( .A1(N144), .A2(N1670), .ZN(N1627) );
  CKND2D0BWPHVT U540 ( .A1(N240), .A2(N1255), .ZN(N1606) );
  CKND0BWPHVT U541 ( .I(N1355), .ZN(N240) );
  CKND2D0BWPHVT U542 ( .A1(N1432), .A2(N1185), .ZN(N1548) );
  AN2D0BWPHVT U543 ( .A1(N13), .A2(N1292), .Z(N1537) );
  CKND0BWPHVT U544 ( .I(N719), .ZN(N1528) );
  CKND2D0BWPHVT U545 ( .A1(N876), .A2(N1132), .ZN(N1523) );
  CKND2D0BWPHVT U546 ( .A1(N1768), .A2(N1366), .ZN(N876) );
  CKND2D0BWPHVT U547 ( .A1(N270), .A2(N1489), .ZN(N1517) );
  CKND2D0BWPHVT U548 ( .A1(N207), .A2(N287), .ZN(N1514) );
  CKND0BWPHVT U549 ( .I(N52), .ZN(N1512) );
  AN2D0BWPHVT U550 ( .A1(N13), .A2(N210), .Z(N150) );
  CKND2D0BWPHVT U551 ( .A1(N12), .A2(N1062), .ZN(N210) );
  CKND2D0BWPHVT U552 ( .A1(N711), .A2(N555), .ZN(N1467) );
  CKND2D0BWPHVT U553 ( .A1(N609), .A2(N513), .ZN(N555) );
  CKND2D0BWPHVT U554 ( .A1(N71), .A2(N266), .ZN(N711) );
  CKND2D0BWPHVT U555 ( .A1(N1235), .A2(N981), .ZN(N1458) );
  CKND0BWPHVT U556 ( .I(N1489), .ZN(N1447) );
  CKND2D0BWPHVT U557 ( .A1(N319), .A2(N2), .ZN(N1443) );
  CKND2D0BWPHVT U558 ( .A1(N923), .A2(N456), .ZN(N1432) );
  CKND2D0BWPHVT U559 ( .A1(N1323), .A2(N1074), .ZN(N1424) );
  CKND2D0BWPHVT U560 ( .A1(N552), .A2(N163), .ZN(N1371) );
  CKND2D0BWPHVT U561 ( .A1(N652), .A2(N1405), .ZN(N137) );
  CKND2D0BWPHVT U562 ( .A1(N897), .A2(N1247), .ZN(N1360) );
  CKND2D0BWPHVT U563 ( .A1(N1036), .A2(N831), .ZN(N897) );
  CKND2D0BWPHVT U564 ( .A1(N334), .A2(N567), .ZN(N1358) );
  CKND2D0BWPHVT U565 ( .A1(N781), .A2(N1502), .ZN(N1355) );
  CKND2D0BWPHVT U566 ( .A1(N1053), .A2(N1048), .ZN(N781) );
  CKND2D0BWPHVT U567 ( .A1(N24), .A2(N528), .ZN(N1344) );
  CKND2D0BWPHVT U568 ( .A1(N449), .A2(N1091), .ZN(N1327) );
  CKND2D0BWPHVT U569 ( .A1(N786), .A2(N320), .ZN(N1292) );
  CKND2D0BWPHVT U570 ( .A1(N523), .A2(N646), .ZN(N320) );
  CKND0BWPHVT U571 ( .I(N290), .ZN(N646) );
  CKND2D0BWPHVT U572 ( .A1(N967), .A2(N290), .ZN(N786) );
  CKND2D0BWPHVT U573 ( .A1(n424), .A2(N149), .ZN(N290) );
  CKND2D0BWPHVT U574 ( .A1(N1452), .A2(N138), .ZN(N1282) );
  CKND2D0BWPHVT U575 ( .A1(N161), .A2(N745), .ZN(N138) );
  CKND2D0BWPHVT U576 ( .A1(N790), .A2(N1136), .ZN(N1452) );
  CKND0BWPHVT U577 ( .I(N302), .ZN(N1255) );
  CKND2D0BWPHVT U578 ( .A1(N683), .A2(N296), .ZN(N302) );
  CKND2D0BWPHVT U579 ( .A1(N1823), .A2(N260), .ZN(N296) );
  CKND0BWPHVT U580 ( .I(N1477), .ZN(N260) );
  CKND2D0BWPHVT U581 ( .A1(N1457), .A2(N1477), .ZN(N683) );
  CKND2D0BWPHVT U582 ( .A1(N1139), .A2(N1569), .ZN(N1477) );
  CKND0BWPHVT U583 ( .I(N1823), .ZN(N1457) );
  CKND2D0BWPHVT U584 ( .A1(N462), .A2(N724), .ZN(N1823) );
  CKND2D0BWPHVT U585 ( .A1(N648), .A2(N1104), .ZN(N1247) );
  CKND0BWPHVT U586 ( .I(N1460), .ZN(N1235) );
  IND2D0BWPHVT U587 ( .A1(N1172), .B1(N1722), .ZN(N1460) );
  CKND2D0BWPHVT U588 ( .A1(N943), .A2(N1326), .ZN(N1233) );
  CKND2D0BWPHVT U589 ( .A1(N406), .A2(N1136), .ZN(N1230) );
  CKND2D0BWPHVT U590 ( .A1(N917), .A2(N1787), .ZN(N1227) );
  CKND2D0BWPHVT U591 ( .A1(N99), .A2(N681), .ZN(N1787) );
  CKND2D0BWPHVT U592 ( .A1(N1408), .A2(N124), .ZN(N917) );
  CKND2D0BWPHVT U593 ( .A1(N1310), .A2(N1575), .ZN(N12) );
  CKND0BWPHVT U594 ( .I(N594), .ZN(N1575) );
  CKND2D0BWPHVT U595 ( .A1(N909), .A2(N227), .ZN(N1185) );
  CKND2D0BWPHVT U596 ( .A1(N919), .A2(N1236), .ZN(N116) );
  CKND2D0BWPHVT U597 ( .A1(N343), .A2(N1577), .ZN(N1236) );
  CKND0BWPHVT U598 ( .I(N977), .ZN(N1577) );
  CKND2D0BWPHVT U599 ( .A1(N386), .A2(N977), .ZN(N919) );
  CKND2D0BWPHVT U600 ( .A1(n424), .A2(N749), .ZN(N977) );
  AN4D0BWPHVT U601 ( .A1(N1204), .A2(N1791), .A3(N77), .A4(N462), .Z(N1156) );
  INR2D0BWPHVT U602 ( .A1(N1176), .B1(N35), .ZN(N1204) );
  AN4D0BWPHVT U603 ( .A1(N1335), .A2(N1364), .A3(n425), .A4(n426), .Z(N1176)
         );
  AN4D0BWPHVT U604 ( .A1(N921), .A2(N376), .A3(N354), .A4(N349), .Z(n426) );
  ND3D0BWPHVT U605 ( .A1(N396), .A2(N1722), .A3(n427), .ZN(N349) );
  ND3D0BWPHVT U606 ( .A1(N1754), .A2(N828), .A3(n428), .ZN(N354) );
  ND3D0BWPHVT U607 ( .A1(N828), .A2(N1189), .A3(n428), .ZN(N376) );
  ND3D0BWPHVT U608 ( .A1(N730), .A2(N253), .A3(n428), .ZN(N921) );
  AN2D0BWPHVT U609 ( .A1(N200), .A2(N1743), .Z(n425) );
  ND3D0BWPHVT U610 ( .A1(N730), .A2(N1633), .A3(n428), .ZN(N1743) );
  AN3D0BWPHVT U611 ( .A1(N243), .A2(N1187), .A3(N396), .Z(n428) );
  ND3D0BWPHVT U612 ( .A1(n427), .A2(N243), .A3(N76), .ZN(N200) );
  NR2D0BWPHVT U613 ( .A1(N543), .A2(N582), .ZN(N76) );
  ND3D0BWPHVT U614 ( .A1(N243), .A2(N1042), .A3(n427), .ZN(N1364) );
  ND3D0BWPHVT U615 ( .A1(n427), .A2(N396), .A3(N694), .ZN(N1335) );
  NR2D0BWPHVT U616 ( .A1(N531), .A2(N591), .ZN(N694) );
  AN3D0BWPHVT U617 ( .A1(N730), .A2(N1187), .A3(N828), .Z(n427) );
  CKND0BWPHVT U618 ( .I(N1330), .ZN(N1187) );
  CKND2D0BWPHVT U619 ( .A1(N1140), .A2(N1052), .ZN(N1137) );
  CKND0BWPHVT U620 ( .I(N1373), .ZN(N1140) );
  XNR2D0BWPHVT U621 ( .A1(N1416), .A2(N1489), .ZN(N1373) );
  CKND2D0BWPHVT U622 ( .A1(n424), .A2(N882), .ZN(N1489) );
  CKND2D0BWPHVT U623 ( .A1(N932), .A2(N1332), .ZN(N1132) );
  CKND2D0BWPHVT U624 ( .A1(N7), .A2(N580), .ZN(N1120) );
  CKND2D0BWPHVT U625 ( .A1(N703), .A2(N802), .ZN(N1093) );
  INR3D0BWPHVT U626 ( .A1(N1791), .B1(N1502), .B2(N77), .ZN(N1088) );
  ND4D0BWPHVT U627 ( .A1(N396), .A2(N828), .A3(N730), .A4(N243), .ZN(N1791) );
  CKND2D0BWPHVT U628 ( .A1(N606), .A2(N222), .ZN(N1073) );
  CKND2D0BWPHVT U629 ( .A1(N766), .A2(N698), .ZN(N222) );
  CKND2D0BWPHVT U630 ( .A1(N438), .A2(N1074), .ZN(N606) );
  CKND2D0BWPHVT U631 ( .A1(N1257), .A2(N594), .ZN(N1062) );
  CKND2D0BWPHVT U632 ( .A1(n424), .A2(N949), .ZN(N594) );
  CKND2D0BWPHVT U633 ( .A1(N755), .A2(N514), .ZN(N1049) );
  CKND2D0BWPHVT U634 ( .A1(N586), .A2(N1501), .ZN(N514) );
  CKND0BWPHVT U635 ( .I(N1096), .ZN(N586) );
  CKND2D0BWPHVT U636 ( .A1(N1096), .A2(N684), .ZN(N755) );
  CKND2D0BWPHVT U637 ( .A1(N4), .A2(N78), .ZN(N1037) );
  AN2D0BWPHVT U638 ( .A1(N13), .A2(N773), .Z(N1025) );
  CKND2D0BWPHVT U639 ( .A1(N722), .A2(N1179), .ZN(N773) );
  CKND2D0BWPHVT U640 ( .A1(N540), .A2(N1383), .ZN(N1179) );
  CKND0BWPHVT U641 ( .I(N1674), .ZN(N1383) );
  CKND0BWPHVT U642 ( .I(N1231), .ZN(N540) );
  CKND2D0BWPHVT U643 ( .A1(N1674), .A2(N1231), .ZN(N722) );
  CKND2D0BWPHVT U644 ( .A1(n424), .A2(N288), .ZN(N1231) );
  NR2D0BWPHVT U645 ( .A1(n429), .A2(N21), .ZN(n424) );
  CKND0BWPHVT U646 ( .I(N35), .ZN(n429) );
  CKND2D0BWPHVT U647 ( .A1(N1020), .A2(N111), .ZN(N35) );
  CKND0BWPHVT U648 ( .I(N724), .ZN(N111) );
  CKND2D0BWPHVT U649 ( .A1(n430), .A2(n431), .ZN(N724) );
  NR4D0BWPHVT U650 ( .A1(N99), .A2(N161), .A3(N660), .A4(N1036), .ZN(n431) );
  CKND0BWPHVT U651 ( .I(N648), .ZN(N1036) );
  ND3D0BWPHVT U652 ( .A1(N8), .A2(n432), .A3(N828), .ZN(N648) );
  CKND0BWPHVT U653 ( .I(N652), .ZN(N660) );
  ND3D0BWPHVT U654 ( .A1(N730), .A2(n432), .A3(N1423), .ZN(N652) );
  CKND0BWPHVT U655 ( .I(N790), .ZN(N161) );
  ND3D0BWPHVT U656 ( .A1(N1633), .A2(n433), .A3(N730), .ZN(N790) );
  CKND0BWPHVT U657 ( .I(N1408), .ZN(N99) );
  ND3D0BWPHVT U658 ( .A1(N1189), .A2(n432), .A3(N253), .ZN(N1408) );
  NR4D0BWPHVT U659 ( .A1(N71), .A2(N26), .A3(N633), .A4(N1683), .ZN(n430) );
  CKND0BWPHVT U660 ( .I(N181), .ZN(N1683) );
  ND3D0BWPHVT U661 ( .A1(n433), .A2(N1189), .A3(N828), .ZN(N181) );
  CKND0BWPHVT U662 ( .I(N319), .ZN(N633) );
  ND3D0BWPHVT U663 ( .A1(N828), .A2(n433), .A3(N1754), .ZN(N319) );
  NR2D0BWPHVT U664 ( .A1(N1100), .A2(N1799), .ZN(N828) );
  CKND0BWPHVT U665 ( .I(N566), .ZN(N26) );
  ND3D0BWPHVT U666 ( .A1(n433), .A2(N253), .A3(N730), .ZN(N566) );
  AN2D0BWPHVT U667 ( .A1(N1722), .A2(n434), .Z(n433) );
  CKND0BWPHVT U668 ( .I(N609), .ZN(N71) );
  ND3D0BWPHVT U669 ( .A1(N253), .A2(n432), .A3(N1754), .ZN(N609) );
  AN2D0BWPHVT U670 ( .A1(N243), .A2(n434), .Z(n432) );
  AN2D0BWPHVT U671 ( .A1(N1042), .A2(N123), .Z(n434) );
  CKND2D0BWPHVT U672 ( .A1(N397), .A2(N1330), .ZN(N123) );
  ND3D0BWPHVT U673 ( .A1(n435), .A2(N1273), .A3(N1824), .ZN(N397) );
  CKND0BWPHVT U674 ( .I(N1139), .ZN(n435) );
  CKND2D0BWPHVT U675 ( .A1(N1502), .A2(N1219), .ZN(N1139) );
  CKND0BWPHVT U676 ( .I(N1048), .ZN(N1219) );
  CKND2D0BWPHVT U677 ( .A1(N1502), .A2(N389), .ZN(N13) );
  CKND0BWPHVT U678 ( .I(N77), .ZN(N389) );
  CKND0BWPHVT U679 ( .I(N1268), .ZN(N1020) );
  CKND2D0BWPHVT U680 ( .A1(N760), .A2(N1711), .ZN(N1018) );
  CKND2D0BWPHVT U681 ( .A1(N165), .A2(N43), .ZN(N1711) );
  CKND0BWPHVT U682 ( .I(N804), .ZN(N43) );
  CKND0BWPHVT U683 ( .I(N23), .ZN(N165) );
  CKND2D0BWPHVT U684 ( .A1(N804), .A2(N23), .ZN(N760) );
  CKND2D0BWPHVT U685 ( .A1(N803), .A2(N1502), .ZN(N23) );
  CKND2D0BWPHVT U686 ( .A1(N1141), .A2(N904), .ZN(N803) );
  CKND2D0BWPHVT U687 ( .A1(N836), .A2(N352), .ZN(N804) );
  CKND2D0BWPHVT U688 ( .A1(N991), .A2(N959), .ZN(N352) );
  CKND0BWPHVT U689 ( .I(N715), .ZN(N959) );
  CKND2D0BWPHVT U690 ( .A1(N715), .A2(N419), .ZN(N836) );
  CKND0BWPHVT U691 ( .I(N991), .ZN(N419) );
  CKND2D0BWPHVT U692 ( .A1(N719), .A2(N1701), .ZN(N991) );
  XNR2D0BWPHVT U693 ( .A1(N602), .A2(N941), .ZN(N719) );
  CKND2D0BWPHVT U694 ( .A1(N1268), .A2(N462), .ZN(N715) );
  ND4D0BWPHVT U695 ( .A1(N1096), .A2(N1172), .A3(n436), .A4(n437), .ZN(N1268)
         );
  NR4D0BWPHVT U696 ( .A1(N1768), .A2(N923), .A3(N552), .A4(N766), .ZN(n437) );
  CKND0BWPHVT U697 ( .I(N438), .ZN(N766) );
  ND3D0BWPHVT U698 ( .A1(N1423), .A2(N730), .A3(n438), .ZN(N438) );
  NR2D0BWPHVT U699 ( .A1(N1682), .A2(N761), .ZN(N730) );
  CKND0BWPHVT U700 ( .I(N449), .ZN(N552) );
  ND4D0BWPHVT U701 ( .A1(n439), .A2(N1633), .A3(N1189), .A4(N243), .ZN(N449)
         );
  NR2D0BWPHVT U702 ( .A1(N1131), .A2(N531), .ZN(N243) );
  CKND0BWPHVT U703 ( .I(N909), .ZN(N923) );
  ND3D0BWPHVT U704 ( .A1(N253), .A2(N1189), .A3(n438), .ZN(N909) );
  CKND0BWPHVT U705 ( .I(N932), .ZN(N1768) );
  ND3D0BWPHVT U706 ( .A1(N1633), .A2(N1189), .A3(n438), .ZN(N932) );
  NR2D0BWPHVT U707 ( .A1(N364), .A2(N1799), .ZN(N1633) );
  NR2D0BWPHVT U708 ( .A1(N323), .A2(N1667), .ZN(n436) );
  CKND0BWPHVT U709 ( .I(N144), .ZN(N1667) );
  CKND2D0BWPHVT U710 ( .A1(n440), .A2(N1754), .ZN(N144) );
  CKND0BWPHVT U711 ( .I(N24), .ZN(N323) );
  ND3D0BWPHVT U712 ( .A1(N1754), .A2(N253), .A3(n438), .ZN(N24) );
  AN3D0BWPHVT U713 ( .A1(N1722), .A2(N1150), .A3(N396), .Z(n438) );
  NR2D0BWPHVT U714 ( .A1(N474), .A2(N543), .ZN(N396) );
  NR2D0BWPHVT U715 ( .A1(N903), .A2(N1682), .ZN(N1754) );
  ND3D0BWPHVT U716 ( .A1(N8), .A2(N253), .A3(n439), .ZN(N1172) );
  NR2D0BWPHVT U717 ( .A1(N569), .A2(N1100), .ZN(N253) );
  NR2D0BWPHVT U718 ( .A1(N224), .A2(N903), .ZN(N8) );
  CKND0BWPHVT U719 ( .I(N761), .ZN(N903) );
  CKND2D0BWPHVT U720 ( .A1(n440), .A2(N1189), .ZN(N1096) );
  NR2D0BWPHVT U721 ( .A1(N224), .A2(N761), .ZN(N1189) );
  CKND2D0BWPHVT U722 ( .A1(N906), .A2(N401), .ZN(N761) );
  CKND2D0BWPHVT U723 ( .A1(N678), .A2(N229), .ZN(N401) );
  CKND2D0BWPHVT U724 ( .A1(N933), .A2(N1536), .ZN(N906) );
  CKND0BWPHVT U725 ( .I(N678), .ZN(N1536) );
  CKND0BWPHVT U726 ( .I(N229), .ZN(N933) );
  CKND2D0BWPHVT U727 ( .A1(N52), .A2(N21), .ZN(N229) );
  CKND2D0BWPHVT U728 ( .A1(N954), .A2(N251), .ZN(N52) );
  CKND2D0BWPHVT U729 ( .A1(N461), .A2(N110), .ZN(N251) );
  CKND2D0BWPHVT U730 ( .A1(N75), .A2(N587), .ZN(N954) );
  CKND0BWPHVT U731 ( .I(N461), .ZN(N587) );
  ND3D0BWPHVT U732 ( .A1(N1134), .A2(N462), .A3(N328), .ZN(N461) );
  CKND0BWPHVT U733 ( .I(N110), .ZN(N75) );
  CKND2D0BWPHVT U734 ( .A1(N763), .A2(N1509), .ZN(N110) );
  CKND2D0BWPHVT U735 ( .A1(N1149), .A2(N471), .ZN(N1509) );
  CKND0BWPHVT U736 ( .I(N1592), .ZN(N471) );
  CKND2D0BWPHVT U737 ( .A1(N1592), .A2(N1016), .ZN(N763) );
  CKND0BWPHVT U738 ( .I(N1149), .ZN(N1016) );
  XNR2D0BWPHVT U739 ( .A1(N1003), .A2(N121), .ZN(N1149) );
  XNR2D0BWPHVT U740 ( .A1(N943), .A2(N1326), .ZN(N1592) );
  CKND0BWPHVT U741 ( .I(N193), .ZN(N943) );
  CKND2D0BWPHVT U742 ( .A1(N992), .A2(N341), .ZN(N193) );
  CKND2D0BWPHVT U743 ( .A1(N416), .A2(N649), .ZN(N341) );
  CKND2D0BWPHVT U744 ( .A1(N1670), .A2(N981), .ZN(N992) );
  CKND0BWPHVT U745 ( .I(N1682), .ZN(N224) );
  CKND2D0BWPHVT U746 ( .A1(N717), .A2(N1518), .ZN(N1682) );
  CKND2D0BWPHVT U747 ( .A1(N873), .A2(N212), .ZN(N1518) );
  CKND0BWPHVT U748 ( .I(N949), .ZN(N212) );
  CKND0BWPHVT U749 ( .I(N1407), .ZN(N873) );
  CKND2D0BWPHVT U750 ( .A1(N949), .A2(N1407), .ZN(N717) );
  CKND2D0BWPHVT U751 ( .A1(N1257), .A2(N21), .ZN(N1407) );
  CKND0BWPHVT U752 ( .I(N1310), .ZN(N1257) );
  XNR2D0BWPHVT U753 ( .A1(N802), .A2(N1113), .ZN(N1310) );
  CKND0BWPHVT U754 ( .I(N703), .ZN(N1113) );
  XNR2D0BWPHVT U755 ( .A1(N4), .A2(N78), .ZN(N703) );
  CKND0BWPHVT U756 ( .I(N207), .ZN(N4) );
  CKND2D0BWPHVT U757 ( .A1(N835), .A2(N379), .ZN(N207) );
  CKND2D0BWPHVT U758 ( .A1(N1104), .A2(N681), .ZN(N379) );
  CKND2D0BWPHVT U759 ( .A1(N124), .A2(N831), .ZN(N835) );
  CKND0BWPHVT U760 ( .I(N496), .ZN(N802) );
  CKND2D0BWPHVT U761 ( .A1(N679), .A2(N1441), .ZN(N496) );
  CKND2D0BWPHVT U762 ( .A1(N973), .A2(N692), .ZN(N1441) );
  CKND0BWPHVT U763 ( .I(N677), .ZN(N692) );
  CKND2D0BWPHVT U764 ( .A1(N677), .A2(N567), .ZN(N679) );
  CKND2D0BWPHVT U765 ( .A1(N1833), .A2(N1242), .ZN(N677) );
  CKND2D0BWPHVT U766 ( .A1(N1465), .A2(N227), .ZN(N1242) );
  CKND0BWPHVT U767 ( .I(N298), .ZN(N1465) );
  CKND2D0BWPHVT U768 ( .A1(N298), .A2(N456), .ZN(N1833) );
  XNR2D0BWPHVT U769 ( .A1(N1095), .A2(N981), .ZN(N298) );
  CKND0BWPHVT U770 ( .I(N1210), .ZN(N1095) );
  ND3D0BWPHVT U771 ( .A1(N462), .A2(N95), .A3(N241), .ZN(N1210) );
  AN3D0BWPHVT U772 ( .A1(N1423), .A2(N1722), .A3(n439), .Z(n440) );
  AN2D0BWPHVT U773 ( .A1(N1042), .A2(N1150), .Z(n439) );
  CKND2D0BWPHVT U774 ( .A1(N537), .A2(N1330), .ZN(N1150) );
  ND3D0BWPHVT U775 ( .A1(N77), .A2(N462), .A3(N1824), .ZN(N1330) );
  IND3D0BWPHVT U776 ( .A1(N1701), .B1(N1273), .B2(N1824), .ZN(N537) );
  CKND2D0BWPHVT U777 ( .A1(N1134), .A2(N1653), .ZN(N1824) );
  CKND2D0BWPHVT U778 ( .A1(N1502), .A2(N148), .ZN(N1701) );
  CKND0BWPHVT U779 ( .I(N904), .ZN(N148) );
  NR2D0BWPHVT U780 ( .A1(N1241), .A2(N474), .ZN(N1042) );
  CKND0BWPHVT U781 ( .I(N582), .ZN(N474) );
  CKND2D0BWPHVT U782 ( .A1(N241), .A2(N1561), .ZN(N582) );
  CKND0BWPHVT U783 ( .I(N543), .ZN(N1241) );
  CKND2D0BWPHVT U784 ( .A1(N1479), .A2(N1195), .ZN(N543) );
  CKND2D0BWPHVT U785 ( .A1(N1775), .A2(N716), .ZN(N1195) );
  CKND0BWPHVT U786 ( .I(N785), .ZN(N716) );
  CKND2D0BWPHVT U787 ( .A1(N288), .A2(N785), .ZN(N1479) );
  CKND2D0BWPHVT U788 ( .A1(N1674), .A2(N21), .ZN(N785) );
  CKND2D0BWPHVT U789 ( .A1(N164), .A2(N1303), .ZN(N1674) );
  CKND2D0BWPHVT U790 ( .A1(N7), .A2(N1569), .ZN(N1303) );
  CKND0BWPHVT U791 ( .I(N580), .ZN(N1569) );
  CKND2D0BWPHVT U792 ( .A1(N1316), .A2(N580), .ZN(N164) );
  CKND2D0BWPHVT U793 ( .A1(N1388), .A2(N1030), .ZN(N580) );
  CKND2D0BWPHVT U794 ( .A1(N64), .A2(N1404), .ZN(N1030) );
  CKND0BWPHVT U795 ( .I(N1440), .ZN(N1404) );
  CKND0BWPHVT U796 ( .I(N1253), .ZN(N64) );
  CKND2D0BWPHVT U797 ( .A1(N1440), .A2(N1253), .ZN(N1388) );
  CKND2D0BWPHVT U798 ( .A1(N90), .A2(N1248), .ZN(N1253) );
  CKND2D0BWPHVT U799 ( .A1(N305), .A2(N899), .ZN(N1248) );
  CKND2D0BWPHVT U800 ( .A1(N1454), .A2(N1431), .ZN(N90) );
  CKND2D0BWPHVT U801 ( .A1(N333), .A2(N1812), .ZN(N1440) );
  CKND2D0BWPHVT U802 ( .A1(N1104), .A2(N745), .ZN(N1812) );
  CKND2D0BWPHVT U803 ( .A1(N1136), .A2(N831), .ZN(N333) );
  CKND0BWPHVT U804 ( .I(N7), .ZN(N1316) );
  XNR2D0BWPHVT U805 ( .A1(N530), .A2(N1511), .ZN(N7) );
  CKND2D0BWPHVT U806 ( .A1(N1053), .A2(N462), .ZN(N1511) );
  XNR2D0BWPHVT U807 ( .A1(N1091), .A2(N1769), .ZN(N530) );
  CKND0BWPHVT U808 ( .I(N1775), .ZN(N288) );
  CKND2D0BWPHVT U809 ( .A1(N1126), .A2(N1561), .ZN(N1775) );
  CKND2D0BWPHVT U810 ( .A1(N95), .A2(N21), .ZN(N1561) );
  NR2D0BWPHVT U811 ( .A1(N1399), .A2(N1131), .ZN(N1722) );
  CKND0BWPHVT U812 ( .I(N591), .ZN(N1131) );
  CKND2D0BWPHVT U813 ( .A1(N767), .A2(N849), .ZN(N591) );
  CKND0BWPHVT U814 ( .I(N531), .ZN(N1399) );
  CKND2D0BWPHVT U815 ( .A1(N268), .A2(N1197), .ZN(N531) );
  CKND2D0BWPHVT U816 ( .A1(N1622), .A2(N538), .ZN(N1197) );
  CKND0BWPHVT U817 ( .I(N749), .ZN(N538) );
  CKND0BWPHVT U818 ( .I(N292), .ZN(N1622) );
  CKND2D0BWPHVT U819 ( .A1(N292), .A2(N749), .ZN(N268) );
  CKND2D0BWPHVT U820 ( .A1(N386), .A2(N21), .ZN(N292) );
  CKND0BWPHVT U821 ( .I(N343), .ZN(N386) );
  XNR2D0BWPHVT U822 ( .A1(N315), .A2(N205), .ZN(N343) );
  CKND2D0BWPHVT U823 ( .A1(N670), .A2(N256), .ZN(N205) );
  CKND2D0BWPHVT U824 ( .A1(N437), .A2(N1166), .ZN(N256) );
  CKND0BWPHVT U825 ( .I(N1328), .ZN(N1166) );
  CKND0BWPHVT U826 ( .I(N1321), .ZN(N437) );
  CKND2D0BWPHVT U827 ( .A1(N1328), .A2(N1321), .ZN(N670) );
  CKND2D0BWPHVT U828 ( .A1(N311), .A2(N1595), .ZN(N1321) );
  CKND2D0BWPHVT U829 ( .A1(N1136), .A2(N1366), .ZN(N1595) );
  CKND2D0BWPHVT U830 ( .A1(N1332), .A2(N745), .ZN(N311) );
  CKND2D0BWPHVT U831 ( .A1(N1141), .A2(N462), .ZN(N1328) );
  CKND0BWPHVT U832 ( .I(N726), .ZN(N315) );
  CKND2D0BWPHVT U833 ( .A1(N258), .A2(N1751), .ZN(N726) );
  CKND2D0BWPHVT U834 ( .A1(N1287), .A2(N441), .ZN(N1751) );
  CKND2D0BWPHVT U835 ( .A1(N1698), .A2(N157), .ZN(N258) );
  CKND0BWPHVT U836 ( .I(N441), .ZN(N157) );
  CKND2D0BWPHVT U837 ( .A1(N276), .A2(N263), .ZN(N441) );
  CKND2D0BWPHVT U838 ( .A1(N1454), .A2(N1769), .ZN(N263) );
  CKND2D0BWPHVT U839 ( .A1(N305), .A2(N1777), .ZN(N276) );
  CKND0BWPHVT U840 ( .I(N1454), .ZN(N305) );
  XNR2D0BWPHVT U841 ( .A1(N1169), .A2(N813), .ZN(N1454) );
  CKND0BWPHVT U842 ( .I(N911), .ZN(N1169) );
  CKND2D0BWPHVT U843 ( .A1(N837), .A2(N1786), .ZN(N911) );
  CKND2D0BWPHVT U844 ( .A1(N2), .A2(N78), .ZN(N1786) );
  CKND0BWPHVT U845 ( .I(N287), .ZN(N78) );
  CKND2D0BWPHVT U846 ( .A1(N287), .A2(N121), .ZN(N837) );
  CKND0BWPHVT U847 ( .I(N2), .ZN(N121) );
  NR2D0BWPHVT U848 ( .A1(N364), .A2(N569), .ZN(N1423) );
  CKND0BWPHVT U849 ( .I(N1799), .ZN(N569) );
  CKND2D0BWPHVT U850 ( .A1(N997), .A2(N1244), .ZN(N1799) );
  CKND2D0BWPHVT U851 ( .A1(N743), .A2(N1029), .ZN(N1244) );
  CKND0BWPHVT U852 ( .I(N882), .ZN(N1029) );
  CKND0BWPHVT U853 ( .I(N1470), .ZN(N743) );
  CKND2D0BWPHVT U854 ( .A1(N1470), .A2(N882), .ZN(N997) );
  CKND2D0BWPHVT U855 ( .A1(N21), .A2(N938), .ZN(N1470) );
  CKND2D0BWPHVT U856 ( .A1(N1312), .A2(N113), .ZN(N938) );
  CKND2D0BWPHVT U857 ( .A1(N270), .A2(N1052), .ZN(N113) );
  CKND0BWPHVT U858 ( .I(N751), .ZN(N1052) );
  CKND0BWPHVT U859 ( .I(N1416), .ZN(N270) );
  CKND2D0BWPHVT U860 ( .A1(N1416), .A2(N751), .ZN(N1312) );
  CKND2D0BWPHVT U861 ( .A1(N1562), .A2(N1238), .ZN(N751) );
  CKND2D0BWPHVT U862 ( .A1(N1763), .A2(N249), .ZN(N1238) );
  CKND0BWPHVT U863 ( .I(N1112), .ZN(N1763) );
  CKND2D0BWPHVT U864 ( .A1(N813), .A2(N1112), .ZN(N1562) );
  ND3D0BWPHVT U865 ( .A1(N462), .A2(N95), .A3(N1126), .ZN(N1112) );
  CKND0BWPHVT U866 ( .I(N1653), .ZN(N95) );
  CKND0BWPHVT U867 ( .I(N249), .ZN(N813) );
  XNR2D0BWPHVT U868 ( .A1(N899), .A2(N941), .ZN(N1416) );
  CKND2D0BWPHVT U869 ( .A1(N593), .A2(N1508), .ZN(N941) );
  CKND2D0BWPHVT U870 ( .A1(N1698), .A2(N1777), .ZN(N1508) );
  CKND0BWPHVT U871 ( .I(N1769), .ZN(N1777) );
  CKND0BWPHVT U872 ( .I(N1287), .ZN(N1698) );
  CKND2D0BWPHVT U873 ( .A1(N1287), .A2(N1769), .ZN(N593) );
  CKND2D0BWPHVT U874 ( .A1(N486), .A2(N1748), .ZN(N1769) );
  CKND2D0BWPHVT U875 ( .A1(N1398), .A2(N1670), .ZN(N1748) );
  CKND2D0BWPHVT U876 ( .A1(N1688), .A2(N649), .ZN(N486) );
  CKND0BWPHVT U877 ( .I(N1398), .ZN(N1688) );
  CKND2D0BWPHVT U878 ( .A1(N562), .A2(N1276), .ZN(N1398) );
  CKND2D0BWPHVT U879 ( .A1(N416), .A2(N1501), .ZN(N1276) );
  CKND2D0BWPHVT U880 ( .A1(N684), .A2(N981), .ZN(N562) );
  CKND0BWPHVT U881 ( .I(N416), .ZN(N981) );
  XNR2D0BWPHVT U882 ( .A1(N1609), .A2(N456), .ZN(N1287) );
  CKND0BWPHVT U883 ( .I(N227), .ZN(N456) );
  CKND0BWPHVT U884 ( .I(N1060), .ZN(N1609) );
  CKND2D0BWPHVT U885 ( .A1(N841), .A2(N1665), .ZN(N1060) );
  CKND2D0BWPHVT U886 ( .A1(N528), .A2(N698), .ZN(N1665) );
  CKND2D0BWPHVT U887 ( .A1(N1074), .A2(N1326), .ZN(N841) );
  CKND0BWPHVT U888 ( .I(N528), .ZN(N1326) );
  CKND0BWPHVT U889 ( .I(N1431), .ZN(N899) );
  CKND2D0BWPHVT U890 ( .A1(N1039), .A2(N1014), .ZN(N1431) );
  CKND2D0BWPHVT U891 ( .A1(N1066), .A2(N124), .ZN(N1039) );
  CKND0BWPHVT U892 ( .I(N1100), .ZN(N364) );
  CKND2D0BWPHVT U893 ( .A1(N812), .A2(N1499), .ZN(N1100) );
  CKND2D0BWPHVT U894 ( .A1(N50), .A2(N149), .ZN(N1499) );
  CKND0BWPHVT U895 ( .I(N271), .ZN(N149) );
  CKND2D0BWPHVT U896 ( .A1(N271), .A2(N1872), .ZN(N812) );
  CKND0BWPHVT U897 ( .I(N50), .ZN(N1872) );
  CKND2D0BWPHVT U898 ( .A1(N967), .A2(N21), .ZN(N50) );
  CKND0BWPHVT U899 ( .I(N523), .ZN(N967) );
  XNR2D0BWPHVT U900 ( .A1(N82), .A2(N481), .ZN(N523) );
  CKND0BWPHVT U901 ( .I(N638), .ZN(N481) );
  XNR2D0BWPHVT U902 ( .A1(N1323), .A2(N698), .ZN(N638) );
  CKND0BWPHVT U903 ( .I(N1074), .ZN(N698) );
  CKND0BWPHVT U904 ( .I(N15), .ZN(N1323) );
  ND3D0BWPHVT U905 ( .A1(N1134), .A2(N462), .A3(N767), .ZN(N15) );
  CKND0BWPHVT U906 ( .I(N1502), .ZN(N462) );
  XNR2D0BWPHVT U907 ( .A1(N567), .A2(N862), .ZN(N82) );
  CKND0BWPHVT U908 ( .I(N334), .ZN(N862) );
  XNR2D0BWPHVT U909 ( .A1(N1142), .A2(N745), .ZN(N334) );
  CKND0BWPHVT U910 ( .I(N1136), .ZN(N745) );
  CKND0BWPHVT U911 ( .I(N406), .ZN(N1142) );
  CKND2D0BWPHVT U912 ( .A1(N187), .A2(N1021), .ZN(N406) );
  CKND2D0BWPHVT U913 ( .A1(N1670), .A2(N777), .ZN(N1021) );
  CKND2D0BWPHVT U914 ( .A1(N1405), .A2(N649), .ZN(N187) );
  CKND0BWPHVT U915 ( .I(N1670), .ZN(N649) );
  CKND0BWPHVT U916 ( .I(N973), .ZN(N567) );
  CKND2D0BWPHVT U917 ( .A1(N92), .A2(N1409), .ZN(N973) );
  CKND2D0BWPHVT U918 ( .A1(N602), .A2(N1501), .ZN(N1409) );
  CKND0BWPHVT U919 ( .I(N684), .ZN(N1501) );
  CKND2D0BWPHVT U920 ( .A1(N650), .A2(N684), .ZN(N92) );
  CKND2D0BWPHVT U921 ( .A1(N328), .A2(N849), .ZN(N271) );
  CKND2D0BWPHVT U922 ( .A1(N1134), .A2(N21), .ZN(N849) );
  CKND0BWPHVT U923 ( .I(N1273), .ZN(N21) );
  CKND2D0BWPHVT U924 ( .A1(N948), .A2(N681), .ZN(N1014) );
  CKND0BWPHVT U925 ( .I(N124), .ZN(N681) );
  CKND0BWPHVT U926 ( .I(N1066), .ZN(N948) );
  CKND2D0BWPHVT U927 ( .A1(N505), .A2(N402), .ZN(N1066) );
  CKND2D0BWPHVT U928 ( .A1(N513), .A2(N777), .ZN(N402) );
  CKND0BWPHVT U929 ( .I(N1405), .ZN(N777) );
  CKND2D0BWPHVT U930 ( .A1(N1405), .A2(N266), .ZN(N505) );
  CKND0BWPHVT U931 ( .I(N1478), .ZN(N1003) );
  CKND2D0BWPHVT U932 ( .A1(N480), .A2(N1565), .ZN(N1478) );
  CKND2D0BWPHVT U933 ( .A1(N513), .A2(N831), .ZN(N1565) );
  CKND0BWPHVT U934 ( .I(N1104), .ZN(N831) );
  CKND2D0BWPHVT U935 ( .A1(N1104), .A2(N266), .ZN(N480) );
  CKND0BWPHVT U936 ( .I(N513), .ZN(N266) );
  CKND0BWPHVT U937 ( .I(N650), .ZN(N602) );
  CKND2D0BWPHVT U938 ( .A1(N969), .A2(N109), .ZN(N650) );
  CKND2D0BWPHVT U939 ( .A1(N1332), .A2(N163), .ZN(N109) );
  CKND0BWPHVT U940 ( .I(N1091), .ZN(N163) );
  CKND2D0BWPHVT U941 ( .A1(N1091), .A2(N1366), .ZN(N969) );
  CKND0BWPHVT U942 ( .I(N1332), .ZN(N1366) );
endmodule

