
module HFC3 (N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670, N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873);

input N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670;
output N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873;
  wire   N906, N1487, N942, N1349, N1744, N1412, N1056, N1320, N888, N1249,
         N1825, N1061, N1723, N467, N2, N77, N124, N227, N249, N287, N416,
         N513, N528, N678, N684, N749, N882, N949, N1074, N1091, N1104, N1134,
         N1136, N1273, N1332, N1405, N1502, N1670, N866, N1272, N17, N251,
         N302, N580, N681, N1648, N555, N1477, N1788, N1372, N461, N582, N1059,
         N745, N615, N698, N397, N652, N541, N740, N553, N477, N1605, N51,
         N245, N1311, N1471, N129, N1146, N529, N757, N423, N647, N1229, N29,
         N546, N1671, N97, N1606, N188, N393, N584, N939, N1573, N970, N471,
         N591, N1419, N1092, N977, N614, N567, N106, N1623, N1708, N116, N1767,
         N156, N234, N405, N1011, N203, N1662, N980, N163, N112, N1870, N381,
         N1051, N549, N668, N692, N297, N271, N1479, N1186, N1303, N885, N945,
         N986, N1310, N117, N714, N1538, N1125, N1789, N402, N209, N788, N131,
         N495, N14, N600, N604, N679, N1546, N1741, N1736, N1548, N1837, N1200,
         N1356, N985, N943, N213, N1393, N298, N1516, N1758, N468, N1574,
         N1547, N1664, N84, N1260, N1600, N551, N1468, N1826, N446, N806, N212,
         N720, N301, N56, N649, N1627, N1351, N1367, N456, N1222, N1759, N687,
         N726, N1773, N1246, N579, N1815, N170, N20, N847, N1208, N1098, N948,
         N576, N777, N1430, N1531, N914, N1279, N1491, N670, N685, N991, N501,
         N815, N1473, N1678, N671, N616, N1131, N1217, N232, N1194, N924,
         N1676, N1427, N1869, N1267, N764, N700, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436;
  assign N164 = N906;
  assign N1435 = N1487;
  assign N833 = N942;
  assign N1255 = N1349;
  assign N81 = N1744;
  assign N323 = N1412;
  assign N427 = N1056;
  assign N325 = N1056;
  assign N564 = N1320;
  assign N1613 = N1320;
  assign N1866 = N888;
  assign N215 = N888;
  assign N178 = N888;
  assign N130 = N888;
  assign N26 = N888;
  assign N1350 = N888;
  assign N1353 = N888;
  assign N765 = N888;
  assign N153 = N1249;
  assign N142 = N1825;
  assign N1015 = N1825;
  assign N602 = N1825;
  assign N974 = N1825;
  assign N1023 = N1825;
  assign N1306 = N1825;
  assign N1301 = N1061;
  assign N1707 = N1723;
  assign N55 = N1723;
  assign N235 = N1723;
  assign N278 = N1723;
  assign N1158 = N467;
  assign N399 = N2;
  assign N1364 = N2;
  assign N878 = N2;
  assign N852 = N2;
  assign N319 = N77;
  assign N99 = N124;
  assign N1342 = N124;
  assign N1127 = N124;
  assign N525 = N124;
  assign N1704 = N227;
  assign N1450 = N227;
  assign N1075 = N227;
  assign N247 = N227;
  assign N1381 = N249;
  assign N1577 = N249;
  assign N770 = N249;
  assign N659 = N249;
  assign N577 = N249;
  assign N101 = N287;
  assign N1872 = N287;
  assign N1509 = N287;
  assign N1 = N287;
  assign N262 = N416;
  assign N1438 = N416;
  assign N1096 = N416;
  assign N1089 = N416;
  assign N531 = N416;
  assign N1190 = N513;
  assign N1404 = N513;
  assign N1386 = N513;
  assign N90 = N513;
  assign N1463 = N528;
  assign N1522 = N528;
  assign N950 = N528;
  assign N669 = N528;
  assign N690 = N678;
  assign N10 = N678;
  assign N1823 = N684;
  assign N1566 = N684;
  assign N1494 = N684;
  assign N1235 = N684;
  assign N113 = N684;
  assign N1277 = N749;
  assign N194 = N749;
  assign N1231 = N882;
  assign N1037 = N882;
  assign N408 = N949;
  assign N177 = N949;
  assign N216 = N1074;
  assign N1775 = N1074;
  assign N1470 = N1074;
  assign N636 = N1074;
  assign N1122 = N1091;
  assign N1798 = N1091;
  assign N1153 = N1091;
  assign N1072 = N1091;
  assign N394 = N1091;
  assign N276 = N1091;
  assign N1757 = N1104;
  assign N794 = N1104;
  assign N620 = N1104;
  assign N35 = N1104;
  assign N1266 = N1134;
  assign N533 = N1134;
  assign N204 = N1136;
  assign N1813 = N1136;
  assign N1309 = N1136;
  assign N1247 = N1136;
  assign N441 = N1136;
  assign N783 = N1273;
  assign N544 = N1273;
  assign N19 = N1332;
  assign N1331 = N1332;
  assign N850 = N1332;
  assign N823 = N1332;
  assign N481 = N1332;
  assign N273 = N1332;
  assign N1111 = N1405;
  assign N1499 = N1405;
  assign N771 = N1405;
  assign N574 = N1405;
  assign N1518 = N1502;
  assign N1497 = N1502;
  assign N1032 = N1502;
  assign N1447 = N1670;
  assign N629 = N1670;
  assign N432 = N1670;
  assign N250 = N1670;
  assign N15 = N1670;
  assign N1274 = N866;
  assign N417 = N866;
  assign N1452 = N1272;
  assign N185 = N1272;
  assign N988 = N17;
  assign N879 = N17;
  assign N293 = N17;
  assign N1534 = N17;
  assign N918 = N251;
  assign N1506 = N302;
  assign N1129 = N302;
  assign N787 = N580;
  assign N1110 = N681;
  assign N360 = N681;
  assign N183 = N1648;
  assign N1174 = N1648;
  assign N1780 = N555;
  assign N1047 = N1477;
  assign N146 = N1477;
  assign N996 = N1477;
  assign N1743 = N1477;
  assign N439 = N1477;
  assign N1838 = N1788;
  assign N1337 = N1372;
  assign N656 = N1372;
  assign N785 = N461;
  assign N1560 = N582;
  assign N429 = N582;
  assign N1012 = N582;
  assign N314 = N1059;
  assign N159 = N745;
  assign N1382 = N615;
  assign N1433 = N698;
  assign N1302 = N698;
  assign N1251 = N698;
  assign N781 = N698;
  assign N752 = N698;
  assign N1237 = N397;
  assign N1033 = N397;
  assign N962 = N397;
  assign N23 = N397;
  assign N496 = N397;
  assign N711 = N652;
  assign N1737 = N541;
  assign N1329 = N541;
  assign N883 = N740;
  assign N96 = N740;
  assign N367 = N740;
  assign N516 = N740;
  assign N1218 = N553;
  assign N1581 = N477;
  assign N1284 = N1605;
  assign N1633 = N51;
  assign N1344 = N51;
  assign N1025 = N51;
  assign N890 = N51;
  assign N1254 = N51;
  assign N1777 = N245;
  assign N1324 = N245;
  assign N644 = N245;
  assign N155 = N245;
  assign N702 = N245;
  assign N308 = N1311;
  assign N1124 = N1311;
  assign N1787 = N1471;
  assign N1774 = N1471;
  assign N1228 = N1471;
  assign N1167 = N1471;
  assign N475 = N1471;
  assign N1685 = N1471;
  assign N857 = N129;
  assign N1058 = N129;
  assign N1856 = N1146;
  assign N1155 = N1146;
  assign N1079 = N1146;
  assign N1071 = N1146;
  assign N1166 = N1146;
  assign N1764 = N529;
  assign N1681 = N757;
  assign N665 = N757;
  assign N867 = N423;
  assign N1183 = N647;
  assign N1117 = N1229;
  assign N539 = N1229;
  assign N378 = N1229;
  assign N284 = N1229;
  assign N148 = N1229;
  assign N733 = N1229;
  assign N1043 = N1229;
  assign N89 = N1229;
  assign N646 = N1229;
  assign N569 = N29;
  assign N1785 = N546;
  assign N1770 = N546;
  assign N484 = N546;
  assign N422 = N546;
  assign N412 = N546;
  assign N182 = N546;
  assign N1388 = N1671;
  assign N1549 = N97;
  assign N1333 = N97;
  assign N1149 = N97;
  assign N372 = N97;
  assign N776 = N97;
  assign N1751 = N1606;
  assign N1373 = N188;
  assign N1026 = N188;
  assign N861 = N188;
  assign N798 = N188;
  assign N1749 = N188;
  assign N1684 = N393;
  assign N1672 = N393;
  assign N759 = N584;
  assign N345 = N584;
  assign N317 = N584;
  assign N187 = N584;
  assign N92 = N584;
  assign N1345 = N584;
  assign N517 = N939;
  assign N494 = N939;
  assign N1696 = N1573;
  assign N5 = N1573;
  assign N1599 = N970;
  assign N1006 = N970;
  assign N1187 = N471;
  assign N1363 = N591;
  assign N98 = N591;
  assign N800 = N1419;
  assign N211 = N1419;
  assign N1556 = N1092;
  assign N275 = N1092;
  assign N1816 = N977;
  assign N1495 = N977;
  assign N1378 = N977;
  assign N1457 = N977;
  assign N1865 = N614;
  assign N1642 = N614;
  assign N1587 = N614;
  assign N1151 = N614;
  assign N1028 = N614;
  assign N639 = N614;
  assign N1602 = N614;
  assign N1532 = N567;
  assign N1638 = N567;
  assign N1409 = N106;
  assign N724 = N106;
  assign N37 = N106;
  assign N827 = N106;
  assign N1178 = N1623;
  assign N1019 = N1623;
  assign N548 = N1708;
  assign N1152 = N1708;
  assign N1423 = N116;
  assign N660 = N116;
  assign N1049 = N1767;
  assign N635 = N156;
  assign N1857 = N234;
  assign N1728 = N405;
  assign N1716 = N405;
  assign N1334 = N405;
  assign N859 = N405;
  assign N1754 = N405;
  assign N1282 = N1011;
  assign N370 = N1011;
  assign N409 = N203;
  assign N1215 = N1662;
  assign N799 = N1662;
  assign N633 = N1662;
  assign N442 = N1662;
  assign N333 = N1662;
  assign N110 = N1662;
  assign N54 = N1662;
  assign N1313 = N1662;
  assign N1140 = N980;
  assign N707 = N980;
  assign N214 = N980;
  assign N851 = N980;
  assign N1198 = N163;
  assign N738 = N163;
  assign N344 = N163;
  assign N645 = N112;
  assign N1008 = N1870;
  assign N755 = N1870;
  assign N479 = N1870;
  assign N340 = N1870;
  assign N169 = N1870;
  assign N946 = N1870;
  assign N63 = N381;
  assign N855 = N1051;
  assign N664 = N549;
  assign N1811 = N668;
  assign N1561 = N692;
  assign N876 = N297;
  assign N457 = N271;
  assign N864 = N1479;
  assign N1384 = N1186;
  assign N510 = N1303;
  assign N274 = N885;
  assign N363 = N945;
  assign N165 = N986;
  assign N1747 = N1310;
  assign N835 = N117;
  assign N1300 = N714;
  assign N438 = N1538;
  assign N920 = N1538;
  assign N121 = N1125;
  assign N1130 = N1789;
  assign N433 = N402;
  assign N627 = N209;
  assign N476 = N788;
  assign N677 = N131;
  assign N1586 = N495;
  assign N1517 = N14;
  assign N1596 = N600;
  assign N352 = N604;
  assign N102 = N679;
  assign N380 = N1546;
  assign N1181 = N1741;
  assign N716 = N1736;
  assign N226 = N1548;
  assign N369 = N1837;
  assign N1214 = N1200;
  assign N594 = N1356;
  assign N192 = N985;
  assign N739 = N943;
  assign N334 = N213;
  assign N1730 = N1393;
  assign N923 = N298;
  assign N1362 = N1516;
  assign N181 = N1758;
  assign N88 = N468;
  assign N1042 = N1574;
  assign N989 = N1547;
  assign N356 = N1547;
  assign N571 = N1547;
  assign N1398 = N1547;
  assign N606 = N1547;
  assign N499 = N1664;
  assign N1480 = N84;
  assign N1210 = N84;
  assign N511 = N1260;
  assign N1385 = N1600;
  assign N195 = N1600;
  assign N421 = N551;
  assign N49 = N1468;
  assign N349 = N1826;
  assign N875 = N1826;
  assign N465 = N446;
  assign N1786 = N806;
  assign N1396 = N806;
  assign N1118 = N212;
  assign N31 = N720;
  assign N512 = N301;
  assign N1540 = N56;
  assign N1064 = N649;
  assign N491 = N649;
  assign N1397 = N1627;
  assign N504 = N1627;
  assign N280 = N1351;
  assign N821 = N1367;
  assign N134 = N456;
  assign N136 = N1222;
  assign N1137 = N1759;
  assign N445 = N687;
  assign N1340 = N687;
  assign N505 = N726;
  assign N1150 = N1773;
  assign N448 = N1246;
  assign N428 = N1246;
  assign N982 = N579;
  assign N1288 = N579;
  assign N898 = N1815;
  assign N834 = N170;
  assign N364 = N20;
  assign N1622 = N847;
  assign N663 = N1208;
  assign N1062 = N1098;
  assign N120 = N948;
  assign N64 = N576;
  assign N122 = N777;
  assign N1276 = N1430;
  assign N1799 = N1531;
  assign N1629 = N914;
  assign N387 = N1279;
  assign N335 = N1491;
  assign N48 = N670;
  assign N266 = N685;
  assign N1808 = N991;
  assign N175 = N501;
  assign N1781 = N815;
  assign N80 = N1473;
  assign N403 = N1678;
  assign N1304 = N671;
  assign N1102 = N671;
  assign N1144 = N671;
  assign N1171 = N616;
  assign N291 = N616;
  assign N1712 = N1131;
  assign N1201 = N1131;
  assign N975 = N1217;
  assign N395 = N1217;
  assign N971 = N232;
  assign N103 = N232;
  assign N1069 = N1194;
  assign N246 = N924;
  assign N1528 = N924;
  assign N128 = N1676;
  assign N655 = N1427;
  assign N1355 = N1869;
  assign N632 = N1267;
  assign N74 = N764;
  assign N38 = N700;

  CKND2D0BWPHVT U470 ( .A1(N582), .A2(N579), .ZN(N997) );
  CKND2D0BWPHVT U471 ( .A1(N671), .A2(N684), .ZN(N991) );
  CKND2D0BWPHVT U472 ( .A1(N1056), .A2(N423), .ZN(N95) );
  CKND2D0BWPHVT U473 ( .A1(N29), .A2(N1870), .ZN(N948) );
  CKND2D0BWPHVT U474 ( .A1(N546), .A2(N990), .ZN(N935) );
  CKND2D0BWPHVT U475 ( .A1(N761), .A2(N1316), .ZN(N880) );
  CKND2D0BWPHVT U476 ( .A1(N796), .A2(N1067), .ZN(N831) );
  CKND2D0BWPHVT U477 ( .A1(N567), .A2(N584), .ZN(N815) );
  CKND2D0BWPHVT U478 ( .A1(N668), .A2(N1670), .ZN(N796) );
  CKND2D0BWPHVT U479 ( .A1(N117), .A2(N287), .ZN(N761) );
  CKND2D0BWPHVT U480 ( .A1(N1573), .A2(N585), .ZN(N760) );
  NR2D0BWPHVT U481 ( .A1(N515), .A2(N1173), .ZN(N728) );
  CKND2D0BWPHVT U482 ( .A1(N912), .A2(N2), .ZN(N723) );
  CKND2D0BWPHVT U483 ( .A1(N78), .A2(N498), .ZN(N697) );
  CKND2D0BWPHVT U484 ( .A1(N271), .A2(N1074), .ZN(N78) );
  CKND2D0BWPHVT U485 ( .A1(N245), .A2(N1229), .ZN(N649) );
  CKND2D0BWPHVT U486 ( .A1(N467), .A2(N1224), .ZN(N617) );
  AN2D0BWPHVT U487 ( .A1(N698), .A2(N1119), .Z(N599) );
  CKND2D0BWPHVT U488 ( .A1(N1338), .A2(N1074), .ZN(N570) );
  CKND2D0BWPHVT U489 ( .A1(N1128), .A2(N1146), .ZN(N543) );
  CKND2D0BWPHVT U490 ( .A1(N286), .A2(N17), .ZN(N535) );
  CKND2D0BWPHVT U491 ( .A1(N140), .A2(N188), .ZN(N534) );
  AN4D0BWPHVT U492 ( .A1(N339), .A2(N454), .A3(N77), .A4(N163), .Z(N515) );
  CKND2D0BWPHVT U493 ( .A1(N981), .A2(N1291), .ZN(N514) );
  CKND2D0BWPHVT U494 ( .A1(N1303), .A2(N1405), .ZN(N981) );
  CKND2D0BWPHVT U495 ( .A1(N795), .A2(N977), .ZN(N498) );
  CKND0BWPHVT U496 ( .I(N271), .ZN(N795) );
  CKND2D0BWPHVT U497 ( .A1(N1825), .A2(N555), .ZN(N495) );
  CKND2D0BWPHVT U498 ( .A1(N1592), .A2(N287), .ZN(N426) );
  CKND2D0BWPHVT U499 ( .A1(N689), .A2(N410), .ZN(N357) );
  CKND2D0BWPHVT U500 ( .A1(N145), .A2(N97), .ZN(N410) );
  CKND2D0BWPHVT U501 ( .A1(N297), .A2(N513), .ZN(N689) );
  INR2D0BWPHVT U502 ( .A1(N1365), .B1(N863), .ZN(N339) );
  CKND2D0BWPHVT U503 ( .A1(N619), .A2(N453), .ZN(N337) );
  CKND2D0BWPHVT U504 ( .A1(N692), .A2(N2), .ZN(N453) );
  CKND2D0BWPHVT U505 ( .A1(N143), .A2(N17), .ZN(N619) );
  CKND2D0BWPHVT U506 ( .A1(N977), .A2(N1406), .ZN(N267) );
  CKND2D0BWPHVT U507 ( .A1(N298), .A2(N1217), .ZN(N213) );
  CKND2D0BWPHVT U508 ( .A1(N180), .A2(N1136), .ZN(N207) );
  CKND2D0BWPHVT U509 ( .A1(N87), .A2(N1720), .ZN(N193) );
  CKND2D0BWPHVT U510 ( .A1(N381), .A2(N416), .ZN(N87) );
  CKND2D0BWPHVT U511 ( .A1(N1200), .A2(N249), .ZN(N1837) );
  CKND2D0BWPHVT U512 ( .A1(N1259), .A2(N1107), .ZN(N1800) );
  AN2D0BWPHVT U513 ( .A1(N698), .A2(N1474), .Z(N1782) );
  CKND2D0BWPHVT U514 ( .A1(N1471), .A2(N1194), .ZN(N1759) );
  CKND2D0BWPHVT U515 ( .A1(N1595), .A2(N546), .ZN(N1720) );
  CKND2D0BWPHVT U516 ( .A1(N444), .A2(N1082), .ZN(N1660) );
  CKND2D0BWPHVT U517 ( .A1(N279), .A2(N1863), .ZN(N444) );
  CKND0BWPHVT U518 ( .I(N230), .ZN(N1863) );
  CKND0BWPHVT U519 ( .I(N22), .ZN(N279) );
  CKND2D0BWPHVT U520 ( .A1(N940), .A2(N419), .ZN(N1641) );
  CKND2D0BWPHVT U521 ( .A1(N1325), .A2(N397), .ZN(N419) );
  CKND2D0BWPHVT U522 ( .A1(N714), .A2(N124), .ZN(N940) );
  CKND2D0BWPHVT U523 ( .A1(N1825), .A2(N888), .ZN(N1627) );
  CKND2D0BWPHVT U524 ( .A1(N756), .A2(N190), .ZN(N1569) );
  CKND2D0BWPHVT U525 ( .A1(N549), .A2(N528), .ZN(N190) );
  CKND2D0BWPHVT U526 ( .A1(N628), .A2(N188), .ZN(N756) );
  CKND2D0BWPHVT U527 ( .A1(N507), .A2(N1779), .ZN(N1562) );
  CKND2D0BWPHVT U528 ( .A1(N972), .A2(N1662), .ZN(N1779) );
  CKND2D0BWPHVT U529 ( .A1(N986), .A2(N1332), .ZN(N507) );
  CKND2D0BWPHVT U530 ( .A1(N745), .A2(N1471), .ZN(N1548) );
  CKND2D0BWPHVT U531 ( .A1(N65), .A2(N1121), .ZN(N1545) );
  CKND2D0BWPHVT U532 ( .A1(N618), .A2(N1471), .ZN(N65) );
  CKND0BWPHVT U533 ( .I(N1479), .ZN(N618) );
  AN2D0BWPHVT U534 ( .A1(N698), .A2(N85), .Z(N1520) );
  CKND2D0BWPHVT U535 ( .A1(N810), .A2(N336), .ZN(N85) );
  CKND2D0BWPHVT U536 ( .A1(N608), .A2(N301), .ZN(N336) );
  CKND2D0BWPHVT U537 ( .A1(N1044), .A2(N911), .ZN(N810) );
  CKND0BWPHVT U538 ( .I(N608), .ZN(N911) );
  CKND2D0BWPHVT U539 ( .A1(n420), .A2(N949), .ZN(N608) );
  CKND2D0BWPHVT U540 ( .A1(N256), .A2(N217), .ZN(N150) );
  CKND2D0BWPHVT U541 ( .A1(N885), .A2(N1091), .ZN(N217) );
  CKND2D0BWPHVT U542 ( .A1(N1544), .A2(N614), .ZN(N256) );
  CKND2D0BWPHVT U543 ( .A1(N1555), .A2(N405), .ZN(N1484) );
  CKND2D0BWPHVT U544 ( .A1(N219), .A2(N1827), .ZN(N1474) );
  CKND2D0BWPHVT U545 ( .A1(N1851), .A2(N547), .ZN(N1827) );
  CKND0BWPHVT U546 ( .I(N901), .ZN(N547) );
  CKND0BWPHVT U547 ( .I(N209), .ZN(N1851) );
  CKND2D0BWPHVT U548 ( .A1(N901), .A2(N209), .ZN(N219) );
  CKND2D0BWPHVT U549 ( .A1(n420), .A2(N749), .ZN(N901) );
  CKND0BWPHVT U550 ( .I(N297), .ZN(N145) );
  CKND2D0BWPHVT U551 ( .A1(N245), .A2(N600), .ZN(N14) );
  CKND2D0BWPHVT U552 ( .A1(N1623), .A2(N1059), .ZN(N1393) );
  CKND0BWPHVT U553 ( .I(N1217), .ZN(N1623) );
  AN2D0BWPHVT U554 ( .A1(N698), .A2(N362), .Z(N1377) );
  CKND2D0BWPHVT U555 ( .A1(N45), .A2(N1336), .ZN(N362) );
  CKND2D0BWPHVT U556 ( .A1(N1568), .A2(N107), .ZN(N45) );
  CKND0BWPHVT U557 ( .I(N1055), .ZN(N1568) );
  CKND2D0BWPHVT U558 ( .A1(N1606), .A2(N51), .ZN(N1367) );
  AN4D0BWPHVT U559 ( .A1(N11), .A2(N1359), .A3(n421), .A4(n422), .Z(N1365) );
  AN4D0BWPHVT U560 ( .A1(N967), .A2(N934), .A3(N440), .A4(N310), .Z(n422) );
  ND3D0BWPHVT U561 ( .A1(n423), .A2(N1428), .A3(N359), .ZN(N310) );
  NR2D0BWPHVT U562 ( .A1(N1356), .A2(N456), .ZN(N359) );
  ND3D0BWPHVT U563 ( .A1(N338), .A2(N478), .A3(n423), .ZN(N440) );
  ND3D0BWPHVT U564 ( .A1(N338), .A2(N392), .A3(n423), .ZN(N934) );
  ND3D0BWPHVT U565 ( .A1(N1428), .A2(N866), .A3(n423), .ZN(N967) );
  AN3D0BWPHVT U566 ( .A1(N791), .A2(N261), .A3(N366), .Z(n423) );
  AN2D0BWPHVT U567 ( .A1(N1807), .A2(N1571), .Z(n421) );
  ND3D0BWPHVT U568 ( .A1(N366), .A2(N1272), .A3(n424), .ZN(N1571) );
  ND3D0BWPHVT U569 ( .A1(N955), .A2(N791), .A3(n424), .ZN(N1807) );
  ND3D0BWPHVT U570 ( .A1(N1675), .A2(N791), .A3(n424), .ZN(N1359) );
  CKND2D0BWPHVT U571 ( .A1(N1491), .A2(N227), .ZN(N1351) );
  CKND2D0BWPHVT U572 ( .A1(N416), .A2(N894), .ZN(N1346) );
  CKND2D0BWPHVT U573 ( .A1(N501), .A2(N1055), .ZN(N1336) );
  AN2D0BWPHVT U574 ( .A1(N698), .A2(N202), .Z(N1318) );
  CKND2D0BWPHVT U575 ( .A1(N805), .A2(N431), .ZN(N202) );
  CKND2D0BWPHVT U576 ( .A1(N129), .A2(N1352), .ZN(N431) );
  CKND0BWPHVT U577 ( .I(N231), .ZN(N1352) );
  CKND2D0BWPHVT U578 ( .A1(N1249), .A2(N231), .ZN(N805) );
  CKND2D0BWPHVT U579 ( .A1(N347), .A2(N1717), .ZN(N231) );
  CKND2D0BWPHVT U580 ( .A1(N84), .A2(N400), .ZN(N1717) );
  CKND2D0BWPHVT U581 ( .A1(N1176), .A2(N1605), .ZN(N347) );
  CKND2D0BWPHVT U582 ( .A1(N1440), .A2(N1146), .ZN(N1316) );
  CKND2D0BWPHVT U583 ( .A1(N930), .A2(N528), .ZN(N13) );
  CKND2D0BWPHVT U584 ( .A1(N666), .A2(N980), .ZN(N1291) );
  CKND2D0BWPHVT U585 ( .A1(N945), .A2(N227), .ZN(N1259) );
  CKND2D0BWPHVT U586 ( .A1(N828), .A2(N252), .ZN(N1230) );
  CKND2D0BWPHVT U587 ( .A1(N21), .A2(N1417), .ZN(N252) );
  CKND2D0BWPHVT U588 ( .A1(N622), .A2(N24), .ZN(N828) );
  CKND0BWPHVT U589 ( .I(N21), .ZN(N24) );
  CKND2D0BWPHVT U590 ( .A1(N485), .A2(N1502), .ZN(N21) );
  CKND2D0BWPHVT U591 ( .A1(N1053), .A2(N1048), .ZN(N485) );
  CKND0BWPHVT U592 ( .I(N1417), .ZN(N622) );
  CKND2D0BWPHVT U593 ( .A1(N846), .A2(N171), .ZN(N1417) );
  CKND2D0BWPHVT U594 ( .A1(N1763), .A2(N811), .ZN(N171) );
  CKND0BWPHVT U595 ( .I(N853), .ZN(N811) );
  CKND2D0BWPHVT U596 ( .A1(N414), .A2(N853), .ZN(N846) );
  CKND2D0BWPHVT U597 ( .A1(N1056), .A2(N480), .ZN(N853) );
  CKND0BWPHVT U598 ( .I(N1763), .ZN(N414) );
  CKND2D0BWPHVT U599 ( .A1(N797), .A2(N163), .ZN(N1763) );
  CKND2D0BWPHVT U600 ( .A1(N1708), .A2(N249), .ZN(N1222) );
  CKND2D0BWPHVT U601 ( .A1(N556), .A2(N12), .ZN(N1212) );
  CKND2D0BWPHVT U602 ( .A1(N1310), .A2(N684), .ZN(N556) );
  CKND2D0BWPHVT U603 ( .A1(N224), .A2(N584), .ZN(N12) );
  CKND0BWPHVT U604 ( .I(N1310), .ZN(N224) );
  CKND2D0BWPHVT U605 ( .A1(N922), .A2(N1256), .ZN(N118) );
  CKND2D0BWPHVT U606 ( .A1(N1051), .A2(N1104), .ZN(N1256) );
  CKND2D0BWPHVT U607 ( .A1(N115), .A2(N106), .ZN(N922) );
  CKND0BWPHVT U608 ( .I(N400), .ZN(N1176) );
  CKND2D0BWPHVT U609 ( .A1(n420), .A2(N882), .ZN(N400) );
  INR3D0BWPHVT U610 ( .A1(N454), .B1(N1502), .B2(N77), .ZN(N1173) );
  ND4D0BWPHVT U611 ( .A1(N338), .A2(N366), .A3(N1428), .A4(N791), .ZN(N454) );
  CKND2D0BWPHVT U612 ( .A1(N1479), .A2(N249), .ZN(N1121) );
  CKND2D0BWPHVT U613 ( .A1(N455), .A2(N191), .ZN(N1119) );
  CKND2D0BWPHVT U614 ( .A1(N964), .A2(N402), .ZN(N191) );
  CKND2D0BWPHVT U615 ( .A1(N1103), .A2(N1791), .ZN(N455) );
  CKND0BWPHVT U616 ( .I(N964), .ZN(N1791) );
  CKND2D0BWPHVT U617 ( .A1(n420), .A2(N678), .ZN(N964) );
  CKND2D0BWPHVT U618 ( .A1(N1554), .A2(N51), .ZN(N1107) );
  CKND0BWPHVT U619 ( .I(N402), .ZN(N1103) );
  ND3D0BWPHVT U620 ( .A1(n424), .A2(N366), .A3(N1376), .ZN(N11) );
  NR2D0BWPHVT U621 ( .A1(N1473), .A2(N679), .ZN(N1376) );
  AN3D0BWPHVT U622 ( .A1(N1428), .A2(N261), .A3(N338), .Z(n424) );
  CKND0BWPHVT U623 ( .I(N9), .ZN(N261) );
  CKND2D0BWPHVT U624 ( .A1(N576), .A2(N1670), .ZN(N1098) );
  CKND2D0BWPHVT U625 ( .A1(N230), .A2(N22), .ZN(N1082) );
  CKND2D0BWPHVT U626 ( .A1(N285), .A2(N1502), .ZN(N22) );
  CKND2D0BWPHVT U627 ( .A1(N1141), .A2(N904), .ZN(N285) );
  CKND2D0BWPHVT U628 ( .A1(N1209), .A2(N1112), .ZN(N230) );
  CKND2D0BWPHVT U629 ( .A1(N1694), .A2(N1070), .ZN(N1112) );
  CKND0BWPHVT U630 ( .I(N1682), .ZN(N1694) );
  CKND2D0BWPHVT U631 ( .A1(N612), .A2(N1682), .ZN(N1209) );
  CKND2D0BWPHVT U632 ( .A1(N1552), .A2(N163), .ZN(N1682) );
  CKND0BWPHVT U633 ( .I(N1070), .ZN(N612) );
  CKND2D0BWPHVT U634 ( .A1(N238), .A2(N858), .ZN(N1070) );
  CKND0BWPHVT U635 ( .I(N653), .ZN(N858) );
  CKND2D0BWPHVT U636 ( .A1(N931), .A2(N502), .ZN(N653) );
  CKND2D0BWPHVT U637 ( .A1(N1320), .A2(N567), .ZN(N502) );
  CKND2D0BWPHVT U638 ( .A1(N1311), .A2(N671), .ZN(N931) );
  CKND0BWPHVT U639 ( .I(N501), .ZN(N107) );
  CKND2D0BWPHVT U640 ( .A1(N686), .A2(N1870), .ZN(N1067) );
  CKND2D0BWPHVT U641 ( .A1(n420), .A2(N757), .ZN(N1055) );
  CKND0BWPHVT U642 ( .I(N301), .ZN(N1044) );
  AN2D0BWPHVT U643 ( .A1(N698), .A2(N651), .Z(N1036) );
  CKND2D0BWPHVT U644 ( .A1(N4), .A2(N149), .ZN(N651) );
  CKND2D0BWPHVT U645 ( .A1(N995), .A2(N906), .ZN(N149) );
  CKND2D0BWPHVT U646 ( .A1(N461), .A2(N1236), .ZN(N4) );
  CKND0BWPHVT U647 ( .I(N995), .ZN(N1236) );
  CKND2D0BWPHVT U648 ( .A1(n420), .A2(N116), .ZN(N995) );
  NR2D0BWPHVT U649 ( .A1(n425), .A2(N203), .ZN(n420) );
  CKND0BWPHVT U650 ( .I(N863), .ZN(n425) );
  CKND2D0BWPHVT U651 ( .A1(N312), .A2(N59), .ZN(N863) );
  CKND0BWPHVT U652 ( .I(N797), .ZN(N59) );
  ND4D0BWPHVT U653 ( .A1(N1479), .A2(N297), .A3(n426), .A4(n427), .ZN(N797) );
  NR4D0BWPHVT U654 ( .A1(N666), .A2(N315), .A3(N1440), .A4(N115), .ZN(n427) );
  CKND0BWPHVT U655 ( .I(N1051), .ZN(N115) );
  ND3D0BWPHVT U656 ( .A1(N1428), .A2(n428), .A3(N184), .ZN(N1051) );
  CKND0BWPHVT U657 ( .I(N117), .ZN(N1440) );
  ND3D0BWPHVT U658 ( .A1(n429), .A2(N1675), .A3(N1428), .ZN(N117) );
  CKND0BWPHVT U659 ( .I(N1303), .ZN(N666) );
  ND3D0BWPHVT U660 ( .A1(N366), .A2(n428), .A3(N109), .ZN(N1303) );
  NR2D0BWPHVT U661 ( .A1(N1325), .A2(N143), .ZN(n426) );
  CKND0BWPHVT U662 ( .I(N692), .ZN(N143) );
  ND3D0BWPHVT U663 ( .A1(N1428), .A2(n429), .A3(N955), .ZN(N692) );
  NR2D0BWPHVT U664 ( .A1(N1600), .A2(N687), .ZN(N1428) );
  CKND0BWPHVT U665 ( .I(N714), .ZN(N1325) );
  ND3D0BWPHVT U666 ( .A1(N1675), .A2(n428), .A3(N392), .ZN(N714) );
  ND3D0BWPHVT U667 ( .A1(N392), .A2(n428), .A3(N955), .ZN(N297) );
  AN3D0BWPHVT U668 ( .A1(N791), .A2(N79), .A3(N866), .Z(n428) );
  ND3D0BWPHVT U669 ( .A1(n429), .A2(N392), .A3(N366), .ZN(N1479) );
  CKND0BWPHVT U670 ( .I(N1552), .ZN(N312) );
  ND4D0BWPHVT U671 ( .A1(N1310), .A2(N271), .A3(n430), .A4(n431), .ZN(N1552)
         );
  NR4D0BWPHVT U672 ( .A1(N972), .A2(N1554), .A3(N1544), .A4(N686), .ZN(n431)
         );
  CKND0BWPHVT U673 ( .I(N668), .ZN(N686) );
  ND3D0BWPHVT U674 ( .A1(N109), .A2(N955), .A3(n432), .ZN(N668) );
  CKND0BWPHVT U675 ( .I(N885), .ZN(N1544) );
  ND4D0BWPHVT U676 ( .A1(N478), .A2(N1675), .A3(n433), .A4(N866), .ZN(N885) );
  AN2D0BWPHVT U677 ( .A1(N1330), .A2(N791), .Z(n433) );
  NR2D0BWPHVT U678 ( .A1(N351), .A2(N679), .ZN(N791) );
  CKND0BWPHVT U679 ( .I(N945), .ZN(N1554) );
  ND3D0BWPHVT U680 ( .A1(N392), .A2(N1675), .A3(n434), .ZN(N945) );
  CKND0BWPHVT U681 ( .I(N986), .ZN(N972) );
  ND3D0BWPHVT U682 ( .A1(N478), .A2(N1675), .A3(n434), .ZN(N986) );
  NR2D0BWPHVT U683 ( .A1(N628), .A2(N1595), .ZN(n430) );
  CKND0BWPHVT U684 ( .I(N381), .ZN(N1595) );
  ND3D0BWPHVT U685 ( .A1(N184), .A2(N392), .A3(n432), .ZN(N381) );
  NR2D0BWPHVT U686 ( .A1(N251), .A2(N652), .ZN(N184) );
  CKND0BWPHVT U687 ( .I(N549), .ZN(N628) );
  ND3D0BWPHVT U688 ( .A1(N955), .A2(N392), .A3(n434), .ZN(N549) );
  NR2D0BWPHVT U689 ( .A1(N553), .A2(N687), .ZN(N392) );
  NR2D0BWPHVT U690 ( .A1(N251), .A2(N806), .ZN(N955) );
  CKND0BWPHVT U691 ( .I(N1538), .ZN(N251) );
  ND3D0BWPHVT U692 ( .A1(N109), .A2(N366), .A3(n434), .ZN(N271) );
  AN3D0BWPHVT U693 ( .A1(N1272), .A2(N1330), .A3(N338), .Z(n434) );
  NR2D0BWPHVT U694 ( .A1(N132), .A2(N1356), .ZN(N338) );
  ND3D0BWPHVT U695 ( .A1(N109), .A2(N1675), .A3(n432), .ZN(N1310) );
  AN3D0BWPHVT U696 ( .A1(N866), .A2(N1330), .A3(N1272), .Z(n432) );
  CKND2D0BWPHVT U697 ( .A1(N9), .A2(N1204), .ZN(N1330) );
  ND3D0BWPHVT U698 ( .A1(N1273), .A2(n435), .A3(N1761), .ZN(N1204) );
  CKND0BWPHVT U699 ( .I(N238), .ZN(n435) );
  CKND2D0BWPHVT U700 ( .A1(N1502), .A2(N1718), .ZN(N238) );
  CKND0BWPHVT U701 ( .I(N904), .ZN(N1718) );
  NR2D0BWPHVT U702 ( .A1(N652), .A2(N1538), .ZN(N1675) );
  CKND0BWPHVT U703 ( .I(N806), .ZN(N652) );
  NR2D0BWPHVT U704 ( .A1(N553), .A2(N529), .ZN(N109) );
  CKND0BWPHVT U705 ( .I(N1600), .ZN(N553) );
  CKND0BWPHVT U706 ( .I(N906), .ZN(N461) );
  CKND2D0BWPHVT U707 ( .A1(N1502), .A2(N615), .ZN(N698) );
  CKND0BWPHVT U708 ( .I(N77), .ZN(N615) );
  CKND2D0BWPHVT U709 ( .A1(N928), .A2(N1812), .ZN(N1014) );
  CKND2D0BWPHVT U710 ( .A1(N1186), .A2(N1136), .ZN(N1812) );
  CKND2D0BWPHVT U711 ( .A1(N315), .A2(N405), .ZN(N928) );
  CKND0BWPHVT U712 ( .I(N1186), .ZN(N315) );
  ND3D0BWPHVT U713 ( .A1(N366), .A2(n429), .A3(N478), .ZN(N1186) );
  NR2D0BWPHVT U714 ( .A1(N529), .A2(N1600), .ZN(N478) );
  CKND2D0BWPHVT U715 ( .A1(N551), .A2(N1468), .ZN(N1600) );
  CKND2D0BWPHVT U716 ( .A1(N477), .A2(N591), .ZN(N1468) );
  CKND0BWPHVT U717 ( .I(N882), .ZN(N591) );
  CKND0BWPHVT U718 ( .I(N1826), .ZN(N477) );
  CKND2D0BWPHVT U719 ( .A1(N1826), .A2(N882), .ZN(N551) );
  CKND2D0BWPHVT U720 ( .A1(N203), .A2(N951), .ZN(N1826) );
  CKND2D0BWPHVT U721 ( .A1(N667), .A2(N1755), .ZN(N951) );
  CKND2D0BWPHVT U722 ( .A1(N129), .A2(N1605), .ZN(N1755) );
  CKND0BWPHVT U723 ( .I(N84), .ZN(N1605) );
  CKND0BWPHVT U724 ( .I(N1249), .ZN(N129) );
  CKND2D0BWPHVT U725 ( .A1(N1249), .A2(N84), .ZN(N667) );
  CKND2D0BWPHVT U726 ( .A1(N446), .A2(N1260), .ZN(N84) );
  CKND2D0BWPHVT U727 ( .A1(N1311), .A2(N1547), .ZN(N1260) );
  CKND0BWPHVT U728 ( .I(N1320), .ZN(N1311) );
  CKND2D0BWPHVT U729 ( .A1(N1320), .A2(N740), .ZN(N446) );
  XNR2D0BWPHVT U730 ( .A1(N1229), .A2(N1825), .ZN(N1320) );
  XNR2D0BWPHVT U731 ( .A1(N1708), .A2(N1471), .ZN(N1249) );
  CKND0BWPHVT U732 ( .I(N1194), .ZN(N1708) );
  ND3D0BWPHVT U733 ( .A1(N163), .A2(N112), .A3(N1126), .ZN(N1194) );
  CKND0BWPHVT U734 ( .I(N687), .ZN(N529) );
  CKND2D0BWPHVT U735 ( .A1(N726), .A2(N1773), .ZN(N687) );
  CKND2D0BWPHVT U736 ( .A1(N1246), .A2(N1487), .ZN(N1773) );
  CKND0BWPHVT U737 ( .I(N939), .ZN(N1487) );
  CKND2D0BWPHVT U738 ( .A1(N939), .A2(N757), .ZN(N726) );
  CKND0BWPHVT U739 ( .I(N1246), .ZN(N757) );
  CKND2D0BWPHVT U740 ( .A1(N328), .A2(N111), .ZN(N1246) );
  CKND2D0BWPHVT U741 ( .A1(N203), .A2(N501), .ZN(N939) );
  CKND2D0BWPHVT U742 ( .A1(N804), .A2(N744), .ZN(N501) );
  CKND2D0BWPHVT U743 ( .A1(N1489), .A2(N30), .ZN(N744) );
  CKND0BWPHVT U744 ( .I(N722), .ZN(N30) );
  CKND2D0BWPHVT U745 ( .A1(N471), .A2(N722), .ZN(N804) );
  CKND2D0BWPHVT U746 ( .A1(N572), .A2(N1090), .ZN(N722) );
  CKND2D0BWPHVT U747 ( .A1(N1767), .A2(N467), .ZN(N1090) );
  CKND2D0BWPHVT U748 ( .A1(N1573), .A2(N371), .ZN(N572) );
  CKND0BWPHVT U749 ( .I(N1767), .ZN(N371) );
  XNR2D0BWPHVT U750 ( .A1(N1555), .A2(N405), .ZN(N1767) );
  CKND0BWPHVT U751 ( .I(N180), .ZN(N1555) );
  CKND2D0BWPHVT U752 ( .A1(N947), .A2(N348), .ZN(N180) );
  CKND2D0BWPHVT U753 ( .A1(N1405), .A2(N1870), .ZN(N348) );
  CKND2D0BWPHVT U754 ( .A1(N1670), .A2(N980), .ZN(N947) );
  CKND0BWPHVT U755 ( .I(N1489), .ZN(N471) );
  XNR2D0BWPHVT U756 ( .A1(N1338), .A2(N977), .ZN(N1489) );
  CKND0BWPHVT U757 ( .I(N1406), .ZN(N1338) );
  ND3D0BWPHVT U758 ( .A1(N1134), .A2(N163), .A3(N767), .ZN(N1406) );
  AN3D0BWPHVT U759 ( .A1(N866), .A2(N79), .A3(N1272), .Z(n429) );
  NR2D0BWPHVT U760 ( .A1(N351), .A2(N580), .ZN(N1272) );
  CKND0BWPHVT U761 ( .I(N679), .ZN(N580) );
  CKND2D0BWPHVT U762 ( .A1(N1741), .A2(N1546), .ZN(N679) );
  CKND2D0BWPHVT U763 ( .A1(N681), .A2(N749), .ZN(N1546) );
  CKND2D0BWPHVT U764 ( .A1(N942), .A2(N970), .ZN(N1741) );
  CKND0BWPHVT U765 ( .I(N749), .ZN(N970) );
  CKND0BWPHVT U766 ( .I(N681), .ZN(N942) );
  CKND2D0BWPHVT U767 ( .A1(N209), .A2(N203), .ZN(N681) );
  CKND2D0BWPHVT U768 ( .A1(N788), .A2(N131), .ZN(N209) );
  CKND2D0BWPHVT U769 ( .A1(N1648), .A2(N924), .ZN(N131) );
  CKND2D0BWPHVT U770 ( .A1(N1061), .A2(N234), .ZN(N788) );
  CKND0BWPHVT U771 ( .I(N924), .ZN(N234) );
  CKND2D0BWPHVT U772 ( .A1(N1676), .A2(N1427), .ZN(N924) );
  CKND2D0BWPHVT U773 ( .A1(N700), .A2(N1869), .ZN(N1427) );
  CKND2D0BWPHVT U774 ( .A1(N156), .A2(N1011), .ZN(N1676) );
  CKND0BWPHVT U775 ( .I(N1869), .ZN(N156) );
  CKND2D0BWPHVT U776 ( .A1(N764), .A2(N1267), .ZN(N1869) );
  CKND2D0BWPHVT U777 ( .A1(N1136), .A2(N1662), .ZN(N1267) );
  CKND2D0BWPHVT U778 ( .A1(N1332), .A2(N405), .ZN(N764) );
  CKND0BWPHVT U779 ( .I(N1648), .ZN(N1061) );
  XNR2D0BWPHVT U780 ( .A1(N555), .A2(N1825), .ZN(N1648) );
  CKND0BWPHVT U781 ( .I(N245), .ZN(N1825) );
  XNR2D0BWPHVT U782 ( .A1(N1606), .A2(N51), .ZN(N245) );
  CKND0BWPHVT U783 ( .I(N1491), .ZN(N1606) );
  CKND2D0BWPHVT U784 ( .A1(N685), .A2(N670), .ZN(N1491) );
  CKND2D0BWPHVT U785 ( .A1(N528), .A2(N977), .ZN(N670) );
  CKND0BWPHVT U786 ( .I(N1074), .ZN(N977) );
  CKND2D0BWPHVT U787 ( .A1(N1074), .A2(N188), .ZN(N685) );
  CKND0BWPHVT U788 ( .I(N600), .ZN(N555) );
  CKND2D0BWPHVT U789 ( .A1(N604), .A2(N1736), .ZN(N600) );
  CKND2D0BWPHVT U790 ( .A1(N1229), .A2(N1477), .ZN(N1736) );
  CKND2D0BWPHVT U791 ( .A1(N888), .A2(N1723), .ZN(N604) );
  CKND0BWPHVT U792 ( .I(N1473), .ZN(N351) );
  CKND2D0BWPHVT U793 ( .A1(N767), .A2(N111), .ZN(N1473) );
  CKND2D0BWPHVT U794 ( .A1(N1134), .A2(N203), .ZN(N111) );
  CKND2D0BWPHVT U795 ( .A1(N9), .A2(N583), .ZN(N79) );
  ND3D0BWPHVT U796 ( .A1(N1273), .A2(n436), .A3(N1761), .ZN(N583) );
  CKND0BWPHVT U797 ( .I(N480), .ZN(n436) );
  CKND2D0BWPHVT U798 ( .A1(N1502), .A2(N1603), .ZN(N480) );
  CKND0BWPHVT U799 ( .I(N1048), .ZN(N1603) );
  ND3D0BWPHVT U800 ( .A1(N77), .A2(N163), .A3(N1761), .ZN(N9) );
  CKND2D0BWPHVT U801 ( .A1(N1134), .A2(N1653), .ZN(N1761) );
  NR2D0BWPHVT U802 ( .A1(N1788), .A2(N132), .ZN(N866) );
  CKND0BWPHVT U803 ( .I(N456), .ZN(N132) );
  CKND2D0BWPHVT U804 ( .A1(N241), .A2(N893), .ZN(N456) );
  CKND0BWPHVT U805 ( .I(N1356), .ZN(N1788) );
  CKND2D0BWPHVT U806 ( .A1(N985), .A2(N943), .ZN(N1356) );
  CKND2D0BWPHVT U807 ( .A1(N232), .A2(N1349), .ZN(N943) );
  CKND0BWPHVT U808 ( .I(N1372), .ZN(N1349) );
  CKND2D0BWPHVT U809 ( .A1(N1372), .A2(N116), .ZN(N985) );
  CKND0BWPHVT U810 ( .I(N232), .ZN(N116) );
  CKND2D0BWPHVT U811 ( .A1(N1126), .A2(N893), .ZN(N232) );
  CKND2D0BWPHVT U812 ( .A1(N112), .A2(N203), .ZN(N893) );
  CKND2D0BWPHVT U813 ( .A1(N906), .A2(N203), .ZN(N1372) );
  CKND2D0BWPHVT U814 ( .A1(N1746), .A2(N162), .ZN(N906) );
  CKND2D0BWPHVT U815 ( .A1(N1056), .A2(N579), .ZN(N162) );
  CKND2D0BWPHVT U816 ( .A1(N582), .A2(N423), .ZN(N1746) );
  CKND0BWPHVT U817 ( .I(N579), .ZN(N423) );
  CKND2D0BWPHVT U818 ( .A1(N1815), .A2(N170), .ZN(N579) );
  CKND2D0BWPHVT U819 ( .A1(N20), .A2(N1678), .ZN(N170) );
  CKND2D0BWPHVT U820 ( .A1(N1092), .A2(N647), .ZN(N1815) );
  CKND0BWPHVT U821 ( .I(N20), .ZN(N647) );
  CKND2D0BWPHVT U822 ( .A1(N847), .A2(N1208), .ZN(N20) );
  CKND2D0BWPHVT U823 ( .A1(N888), .A2(N614), .ZN(N1208) );
  CKND0BWPHVT U824 ( .I(N1229), .ZN(N888) );
  CKND2D0BWPHVT U825 ( .A1(N1229), .A2(N1091), .ZN(N847) );
  XNR2D0BWPHVT U826 ( .A1(N29), .A2(N1870), .ZN(N1229) );
  CKND0BWPHVT U827 ( .I(N576), .ZN(N29) );
  CKND2D0BWPHVT U828 ( .A1(N777), .A2(N1430), .ZN(N576) );
  CKND2D0BWPHVT U829 ( .A1(N684), .A2(N546), .ZN(N1430) );
  CKND2D0BWPHVT U830 ( .A1(N416), .A2(N584), .ZN(N777) );
  CKND0BWPHVT U831 ( .I(N1678), .ZN(N1092) );
  CKND2D0BWPHVT U832 ( .A1(N1053), .A2(N163), .ZN(N1678) );
  CKND0BWPHVT U833 ( .I(N1056), .ZN(N582) );
  XNR2D0BWPHVT U834 ( .A1(N1059), .A2(N1217), .ZN(N1056) );
  CKND2D0BWPHVT U835 ( .A1(N921), .A2(N1192), .ZN(N1217) );
  CKND2D0BWPHVT U836 ( .A1(N1104), .A2(N405), .ZN(N1192) );
  CKND0BWPHVT U837 ( .I(N1136), .ZN(N405) );
  CKND2D0BWPHVT U838 ( .A1(N1136), .A2(N106), .ZN(N921) );
  CKND0BWPHVT U839 ( .I(N298), .ZN(N1059) );
  CKND2D0BWPHVT U840 ( .A1(N1758), .A2(N1516), .ZN(N298) );
  CKND2D0BWPHVT U841 ( .A1(N1477), .A2(N1547), .ZN(N1516) );
  CKND2D0BWPHVT U842 ( .A1(N1723), .A2(N740), .ZN(N1758) );
  CKND0BWPHVT U843 ( .I(N1547), .ZN(N740) );
  CKND2D0BWPHVT U844 ( .A1(N56), .A2(N1664), .ZN(N1547) );
  CKND2D0BWPHVT U845 ( .A1(N1531), .A2(N124), .ZN(N1664) );
  CKND2D0BWPHVT U846 ( .A1(N1671), .A2(N397), .ZN(N56) );
  CKND0BWPHVT U847 ( .I(N1531), .ZN(N1671) );
  CKND2D0BWPHVT U848 ( .A1(N914), .A2(N1279), .ZN(N1531) );
  CKND2D0BWPHVT U849 ( .A1(N1405), .A2(N97), .ZN(N1279) );
  CKND2D0BWPHVT U850 ( .A1(N513), .A2(N980), .ZN(N914) );
  CKND0BWPHVT U851 ( .I(N1405), .ZN(N980) );
  CKND0BWPHVT U852 ( .I(N1477), .ZN(N1723) );
  XNR2D0BWPHVT U853 ( .A1(N745), .A2(N1471), .ZN(N1477) );
  CKND0BWPHVT U854 ( .I(N249), .ZN(N1471) );
  CKND0BWPHVT U855 ( .I(N1200), .ZN(N745) );
  CKND2D0BWPHVT U856 ( .A1(N468), .A2(N1574), .ZN(N1200) );
  CKND2D0BWPHVT U857 ( .A1(N287), .A2(N17), .ZN(N1574) );
  CKND2D0BWPHVT U858 ( .A1(N2), .A2(N1146), .ZN(N468) );
  NR2D0BWPHVT U859 ( .A1(N1538), .A2(N806), .ZN(N366) );
  CKND2D0BWPHVT U860 ( .A1(N720), .A2(N212), .ZN(N806) );
  CKND2D0BWPHVT U861 ( .A1(N1744), .A2(N1419), .ZN(N212) );
  CKND0BWPHVT U862 ( .I(N949), .ZN(N1419) );
  CKND0BWPHVT U863 ( .I(N541), .ZN(N1744) );
  CKND2D0BWPHVT U864 ( .A1(N541), .A2(N949), .ZN(N720) );
  CKND2D0BWPHVT U865 ( .A1(N203), .A2(N301), .ZN(N541) );
  CKND2D0BWPHVT U866 ( .A1(N1391), .A2(N1248), .ZN(N301) );
  CKND2D0BWPHVT U867 ( .A1(N536), .A2(N1842), .ZN(N1248) );
  CKND0BWPHVT U868 ( .I(N384), .ZN(N1842) );
  CKND0BWPHVT U869 ( .I(N42), .ZN(N536) );
  CKND2D0BWPHVT U870 ( .A1(N42), .A2(N384), .ZN(N1391) );
  XNR2D0BWPHVT U871 ( .A1(N1128), .A2(N1146), .ZN(N384) );
  CKND0BWPHVT U872 ( .I(N287), .ZN(N1146) );
  CKND0BWPHVT U873 ( .I(N1592), .ZN(N1128) );
  CKND2D0BWPHVT U874 ( .A1(N425), .A2(N1244), .ZN(N1592) );
  CKND2D0BWPHVT U875 ( .A1(N124), .A2(N106), .ZN(N1244) );
  CKND2D0BWPHVT U876 ( .A1(N1104), .A2(N397), .ZN(N425) );
  CKND0BWPHVT U877 ( .I(N124), .ZN(N397) );
  XNR2D0BWPHVT U878 ( .A1(N585), .A2(N467), .ZN(N42) );
  CKND0BWPHVT U879 ( .I(N1573), .ZN(N467) );
  XNR2D0BWPHVT U880 ( .A1(N567), .A2(N584), .ZN(N1573) );
  CKND0BWPHVT U881 ( .I(N684), .ZN(N584) );
  CKND0BWPHVT U882 ( .I(N671), .ZN(N567) );
  CKND2D0BWPHVT U883 ( .A1(N616), .A2(N1131), .ZN(N671) );
  CKND2D0BWPHVT U884 ( .A1(N1332), .A2(N614), .ZN(N1131) );
  CKND0BWPHVT U885 ( .I(N1091), .ZN(N614) );
  CKND2D0BWPHVT U886 ( .A1(N1091), .A2(N1662), .ZN(N616) );
  CKND0BWPHVT U887 ( .I(N1332), .ZN(N1662) );
  CKND0BWPHVT U888 ( .I(N1224), .ZN(N585) );
  CKND2D0BWPHVT U889 ( .A1(N8), .A2(N346), .ZN(N1224) );
  CKND2D0BWPHVT U890 ( .A1(N1523), .A2(N51), .ZN(N346) );
  CKND0BWPHVT U891 ( .I(N227), .ZN(N51) );
  CKND2D0BWPHVT U892 ( .A1(N809), .A2(N227), .ZN(N8) );
  CKND0BWPHVT U893 ( .I(N1523), .ZN(N809) );
  XNR2D0BWPHVT U894 ( .A1(N894), .A2(N546), .ZN(N1523) );
  CKND0BWPHVT U895 ( .I(N990), .ZN(N894) );
  ND3D0BWPHVT U896 ( .A1(N163), .A2(N112), .A3(N241), .ZN(N990) );
  CKND0BWPHVT U897 ( .I(N1653), .ZN(N112) );
  CKND2D0BWPHVT U898 ( .A1(N1789), .A2(N1125), .ZN(N1538) );
  CKND2D0BWPHVT U899 ( .A1(N1412), .A2(N393), .ZN(N1125) );
  CKND0BWPHVT U900 ( .I(N678), .ZN(N393) );
  CKND0BWPHVT U901 ( .I(N302), .ZN(N1412) );
  CKND2D0BWPHVT U902 ( .A1(N302), .A2(N678), .ZN(N1789) );
  CKND2D0BWPHVT U903 ( .A1(N203), .A2(N402), .ZN(N302) );
  CKND2D0BWPHVT U904 ( .A1(N648), .A2(N1219), .ZN(N402) );
  CKND2D0BWPHVT U905 ( .A1(N469), .A2(N958), .ZN(N1219) );
  CKND0BWPHVT U906 ( .I(N487), .ZN(N958) );
  CKND0BWPHVT U907 ( .I(N1714), .ZN(N469) );
  CKND2D0BWPHVT U908 ( .A1(N487), .A2(N1714), .ZN(N648) );
  CKND2D0BWPHVT U909 ( .A1(N375), .A2(N32), .ZN(N1714) );
  CKND2D0BWPHVT U910 ( .A1(N897), .A2(N390), .ZN(N32) );
  CKND0BWPHVT U911 ( .I(N377), .ZN(N390) );
  CKND2D0BWPHVT U912 ( .A1(N377), .A2(N277), .ZN(N375) );
  CKND0BWPHVT U913 ( .I(N897), .ZN(N277) );
  XNR2D0BWPHVT U914 ( .A1(N140), .A2(N188), .ZN(N897) );
  CKND0BWPHVT U915 ( .I(N528), .ZN(N188) );
  CKND0BWPHVT U916 ( .I(N930), .ZN(N140) );
  CKND2D0BWPHVT U917 ( .A1(N1792), .A2(N1197), .ZN(N930) );
  CKND2D0BWPHVT U918 ( .A1(N1670), .A2(N546), .ZN(N1197) );
  CKND0BWPHVT U919 ( .I(N416), .ZN(N546) );
  CKND2D0BWPHVT U920 ( .A1(N416), .A2(N1870), .ZN(N1792) );
  CKND0BWPHVT U921 ( .I(N1670), .ZN(N1870) );
  XNR2D0BWPHVT U922 ( .A1(N286), .A2(N17), .ZN(N377) );
  CKND0BWPHVT U923 ( .I(N2), .ZN(N17) );
  CKND0BWPHVT U924 ( .I(N912), .ZN(N286) );
  CKND2D0BWPHVT U925 ( .A1(N839), .A2(N789), .ZN(N912) );
  CKND2D0BWPHVT U926 ( .A1(N1104), .A2(N97), .ZN(N789) );
  CKND0BWPHVT U927 ( .I(N513), .ZN(N97) );
  CKND2D0BWPHVT U928 ( .A1(N513), .A2(N106), .ZN(N839) );
  CKND0BWPHVT U929 ( .I(N1104), .ZN(N106) );
  ND3D0BWPHVT U930 ( .A1(N1134), .A2(N163), .A3(N328), .ZN(N487) );
  CKND0BWPHVT U931 ( .I(N1273), .ZN(N203) );
  CKND0BWPHVT U932 ( .I(N700), .ZN(N1011) );
  CKND2D0BWPHVT U933 ( .A1(N1141), .A2(N163), .ZN(N700) );
  CKND0BWPHVT U934 ( .I(N1502), .ZN(N163) );
endmodule

