
module Circuit (N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670, N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873);

input N2, N77, N124, N227, N241, N249, N287, N328, N416, N513, N528, N678, N684, N749, N767, N882, N904, N949, N1048, N1053, N1074, N1091, N1104, N1126, N1134, N1136, N1141, N1273, N1332, N1405, N1502, N1653, N1670;
output N47, N208, N233, N385, N411, N472, N643, N854, N963, N978, N999, N1108, N1109, N1143, N1206, N1211, N1305, N1368, N1486, N1590, N1597, N1615, N1731, N1855, N1873;
  wire   N638, N1097, N299, N1801, N964, N112, N1407, N945, N309, N1297, N1828,
         N909, N1317, N1677, N1760, N2, N77, N124, N227, N249, N287, N416,
         N513, N528, N678, N684, N749, N882, N949, N1074, N1091, N1104, N1134,
         N1136, N1273, N1332, N1405, N1502, N1670, N374, N1802, N509, N1319,
         N1324, N240, N1783, N1383, N1369, N1139, N1018, N357, N628, N108,
         N1252, N1803, N127, N442, N21, N1439, N30, N1806, N1307, N368, N93,
         N805, N648, N316, N1559, N947, N187, N218, N1265, N928, N1525, N1078,
         N1521, N231, N1000, N206, N868, N456, N338, N1666, N876, N1658, N1441,
         N1414, N1449, N1432, N1693, N590, N1604, N1343, N290, N340, N151,
         N490, N1840, N502, N526, N779, N745, N29, N1035, N480, N75, N1073,
         N428, N708, N1236, N1588, N1352, N973, N898, N1168, N153, N673, N298,
         N110, N242, N1189, N1101, N1213, N1422, N1444, N736, N1, N1208, N1745,
         N440, N1613, N966, N825, N1207, N361, N1500, N1645, N1709, N1692,
         N1183, N730, N78, N663, N687, N1360, N1729, N1221, N841, N1393, N1591,
         N1415, N1009, N1700, N1434, N1389, N581, N89, N1830, N596, N465,
         N1589, N1162, N1261, N1185, N235, N1046, N790, N707, N1130, N1356,
         N1437, N1541, N1861, N661, N746, N1069, N1527, N1039, N239, N1298,
         N907, N1462, N1253, N633, N786, N642, N1425, N458, N1245, N1834, N258,
         N727, N974, N1619, N1835, N156, N543, N1117, N48, N1536, N397, N1579,
         N297, N1466, N33, N1794, N146, N984, N753, N1164, N1836, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435;
  assign N447 = N638;
  assign N1481 = N1097;
  assign N372 = N1097;
  assign N574 = N1097;
  assign N524 = N1097;
  assign N1868 = N299;
  assign N322 = N299;
  assign N19 = N1801;
  assign N248 = N964;
  assign N87 = N112;
  assign N467 = N1407;
  assign N1535 = N945;
  assign N895 = N945;
  assign N763 = N945;
  assign N292 = N945;
  assign N271 = N945;
  assign N56 = N945;
  assign N1308 = N945;
  assign N50 = N945;
  assign N1458 = N309;
  assign N698 = N1297;
  assign N283 = N1828;
  assign N423 = N909;
  assign N53 = N909;
  assign N1311 = N909;
  assign N757 = N909;
  assign N535 = N1317;
  assign N1443 = N1317;
  assign N193 = N1317;
  assign N548 = N1317;
  assign N656 = N1317;
  assign N748 = N1317;
  assign N1251 = N1677;
  assign N1116 = N1760;
  assign N1184 = N2;
  assign N1199 = N2;
  assign N1094 = N2;
  assign N137 = N2;
  assign N344 = N77;
  assign N289 = N124;
  assign N729 = N124;
  assign N304 = N124;
  assign N114 = N124;
  assign N229 = N227;
  assign N1287 = N227;
  assign N773 = N227;
  assign N518 = N227;
  assign N1392 = N249;
  assign N1191 = N249;
  assign N717 = N249;
  assign N255 = N249;
  assign N209 = N249;
  assign N497 = N287;
  assign N1329 = N287;
  assign N1157 = N287;
  assign N710 = N287;
  assign N561 = N416;
  assign N768 = N416;
  assign N333 = N416;
  assign N168 = N416;
  assign N105 = N416;
  assign N1611 = N513;
  assign N1656 = N513;
  assign N1120 = N513;
  assign N1059 = N513;
  assign N150 = N528;
  assign N1483 = N528;
  assign N775 = N528;
  assign N173 = N528;
  assign N96 = N678;
  assign N54 = N678;
  assign N1179 = N684;
  assign N1776 = N684;
  assign N1558 = N684;
  assign N670 = N684;
  assign N260 = N684;
  assign N1375 = N749;
  assign N514 = N749;
  assign N715 = N882;
  assign N406 = N882;
  assign N544 = N949;
  assign N487 = N949;
  assign N766 = N1074;
  assign N877 = N1074;
  assign N370 = N1074;
  assign N141 = N1074;
  assign N1687 = N1091;
  assign N1400 = N1091;
  assign N1217 = N1091;
  assign N851 = N1091;
  assign N655 = N1091;
  assign N88 = N1091;
  assign N1100 = N1104;
  assign N1673 = N1104;
  assign N1427 = N1104;
  assign N1295 = N1104;
  assign N336 = N1134;
  assign N41 = N1134;
  assign N107 = N1136;
  assign N1281 = N1136;
  assign N728 = N1136;
  assign N672 = N1136;
  assign N403 = N1136;
  assign N1275 = N1273;
  assign N523 = N1273;
  assign N1543 = N1332;
  assign N1601 = N1332;
  assign N1271 = N1332;
  assign N1024 = N1332;
  assign N784 = N1332;
  assign N335 = N1332;
  assign N1814 = N1405;
  assign N1420 = N1405;
  assign N878 = N1405;
  assign N280 = N1405;
  assign N1690 = N1502;
  assign N1030 = N1502;
  assign N323 = N1502;
  assign N459 = N1670;
  assign N1564 = N1670;
  assign N1544 = N1670;
  assign N1081 = N1670;
  assign N471 = N1670;
  assign N799 = N374;
  assign N721 = N374;
  assign N1635 = N1802;
  assign N522 = N1802;
  assign N1533 = N509;
  assign N777 = N509;
  assign N444 = N509;
  assign N609 = N509;
  assign N1387 = N1319;
  assign N282 = N1319;
  assign N220 = N1324;
  assign N376 = N240;
  assign N1732 = N1783;
  assign N910 = N1783;
  assign N880 = N1383;
  assign N1793 = N1369;
  assign N1411 = N1369;
  assign N1313 = N1139;
  assign N599 = N1018;
  assign N379 = N1018;
  assign N1639 = N357;
  assign N621 = N628;
  assign N623 = N628;
  assign N1222 = N108;
  assign N1557 = N1252;
  assign N189 = N1252;
  assign N1351 = N1252;
  assign N92 = N1252;
  assign N147 = N1252;
  assign N1228 = N1803;
  assign N756 = N127;
  assign N1854 = N442;
  assign N1403 = N442;
  assign N1335 = N442;
  assign N1175 = N442;
  assign N1106 = N442;
  assign N1782 = N21;
  assign N1290 = N21;
  assign N1289 = N21;
  assign N846 = N21;
  assign N1103 = N21;
  assign N1076 = N1439;
  assign N154 = N30;
  assign N1829 = N1806;
  assign N1057 = N1806;
  assign N1702 = N1307;
  assign N451 = N1307;
  assign N693 = N1307;
  assign N965 = N1307;
  assign N486 = N1307;
  assign N874 = N368;
  assign N1864 = N93;
  assign N713 = N805;
  assign N86 = N805;
  assign N1372 = N648;
  assign N1083 = N648;
  assign N484 = N648;
  assign N274 = N648;
  assign N1739 = N648;
  assign N1631 = N316;
  assign N1680 = N316;
  assign N892 = N1559;
  assign N669 = N1559;
  assign N68 = N1559;
  assign N836 = N1559;
  assign N1019 = N1559;
  assign N264 = N947;
  assign N1733 = N187;
  assign N674 = N187;
  assign N351 = N187;
  assign N326 = N187;
  assign N238 = N187;
  assign N473 = N187;
  assign N941 = N218;
  assign N818 = N218;
  assign N396 = N218;
  assign N130 = N218;
  assign N222 = N218;
  assign N785 = N1265;
  assign N1087 = N1265;
  assign N192 = N928;
  assign N625 = N1525;
  assign N1734 = N1078;
  assign N1573 = N1521;
  assign N1482 = N1521;
  assign N665 = N1521;
  assign N637 = N1521;
  assign N433 = N1521;
  assign N3 = N1521;
  assign N1695 = N1521;
  assign N510 = N1521;
  assign N998 = N1521;
  assign N499 = N231;
  assign N1831 = N1000;
  assign N906 = N1000;
  assign N732 = N1000;
  assign N493 = N1000;
  assign N140 = N1000;
  assign N1293 = N1000;
  assign N1399 = N206;
  assign N1797 = N868;
  assign N742 = N868;
  assign N626 = N868;
  assign N594 = N868;
  assign N1539 = N868;
  assign N527 = N456;
  assign N1874 = N338;
  assign N1566 = N338;
  assign N1285 = N338;
  assign N195 = N338;
  assign N118 = N338;
  assign N983 = N1666;
  assign N232 = N1666;
  assign N1524 = N876;
  assign N1410 = N876;
  assign N525 = N876;
  assign N265 = N876;
  assign N139 = N876;
  assign N960 = N876;
  assign N1232 = N1658;
  assign N1832 = N1441;
  assign N199 = N1441;
  assign N1058 = N1414;
  assign N1254 = N1449;
  assign N601 = N1449;
  assign N391 = N1432;
  assign N1381 = N1693;
  assign N556 = N1693;
  assign N1691 = N590;
  assign N1621 = N590;
  assign N45 = N1604;
  assign N404 = N1604;
  assign N389 = N1343;
  assign N136 = N1343;
  assign N81 = N1343;
  assign N12 = N1343;
  assign N161 = N290;
  assign N1361 = N290;
  assign N948 = N340;
  assign N454 = N340;
  assign N267 = N340;
  assign N157 = N340;
  assign N80 = N340;
  assign N62 = N340;
  assign N1029 = N340;
  assign N1027 = N151;
  assign N348 = N151;
  assign N16 = N151;
  assign N4 = N151;
  assign N1778 = N490;
  assign N582 = N490;
  assign N843 = N1840;
  assign N1192 = N1840;
  assign N838 = N502;
  assign N776 = N502;
  assign N144 = N526;
  assign N1082 = N779;
  assign N654 = N745;
  assign N1649 = N29;
  assign N1363 = N29;
  assign N545 = N29;
  assign N286 = N29;
  assign N937 = N29;
  assign N1186 = N1035;
  assign N930 = N1035;
  assign N1659 = N480;
  assign N1779 = N75;
  assign N1668 = N75;
  assign N1582 = N75;
  assign N1260 = N75;
  assign N469 = N75;
  assign N445 = N75;
  assign N343 = N75;
  assign N1657 = N75;
  assign N1726 = N1073;
  assign N1259 = N1073;
  assign N353 = N1073;
  assign N1719 = N1073;
  assign N1738 = N428;
  assign N1365 = N428;
  assign N587 = N428;
  assign N1839 = N708;
  assign N1195 = N1236;
  assign N816 = N1236;
  assign N630 = N1236;
  assign N201 = N1236;
  assign N183 = N1236;
  assign N1137 = N1236;
  assign N418 = N1588;
  assign N1581 = N1352;
  assign N1135 = N973;
  assign N1358 = N898;
  assign N325 = N1168;
  assign N1270 = N153;
  assign N1594 = N673;
  assign N492 = N298;
  assign N520 = N110;
  assign N1431 = N242;
  assign N562 = N1189;
  assign N1147 = N1101;
  assign N82 = N1213;
  assign N101 = N1422;
  assign N758 = N1444;
  assign N402 = N736;
  assign N237 = N1;
  assign N126 = N1;
  assign N377 = N1208;
  assign N739 = N1745;
  assign N866 = N440;
  assign N26 = N1613;
  assign N288 = N966;
  assign N1844 = N825;
  assign N1650 = N1207;
  assign N1721 = N361;
  assign N1740 = N1500;
  assign N275 = N1645;
  assign N35 = N1709;
  assign N1250 = N1692;
  assign N857 = N1183;
  assign N395 = N730;
  assign N245 = N78;
  assign N165 = N663;
  assign N552 = N687;
  assign N1550 = N1360;
  assign N200 = N1729;
  assign N1016 = N1221;
  assign N1618 = N841;
  assign N1660 = N841;
  assign N792 = N841;
  assign N1647 = N1393;
  assign N302 = N1591;
  assign N5 = N1415;
  assign N252 = N1009;
  assign N774 = N1700;
  assign N537 = N1434;
  assign N1051 = N1389;
  assign N450 = N581;
  assign N1475 = N581;
  assign N117 = N89;
  assign N624 = N1830;
  assign N1771 = N596;
  assign N226 = N596;
  assign N1380 = N465;
  assign N682 = N1589;
  assign N1753 = N1589;
  assign N462 = N1162;
  assign N796 = N1261;
  assign N1578 = N1185;
  assign N143 = N235;
  assign N571 = N235;
  assign N607 = N1046;
  assign N470 = N1046;
  assign N1429 = N790;
  assign N1624 = N707;
  assign N987 = N1130;
  assign N1334 = N1356;
  assign N312 = N1356;
  assign N554 = N1437;
  assign N1284 = N1541;
  assign N806 = N1861;
  assign N315 = N1861;
  assign N133 = N661;
  assign N123 = N746;
  assign N61 = N1069;
  assign N916 = N1069;
  assign N17 = N1527;
  assign N1426 = N1527;
  assign N1348 = N1039;
  assign N46 = N239;
  assign N178 = N1298;
  assign N1336 = N907;
  assign N1145 = N1462;
  assign N542 = N1253;
  assign N1860 = N633;
  assign N1099 = N786;
  assign N1551 = N642;
  assign N1262 = N1425;
  assign N84 = N458;
  assign N622 = N1245;
  assign N1005 = N1834;
  assign N463 = N258;
  assign N1725 = N727;
  assign N215 = N974;
  assign N1593 = N1619;
  assign N1153 = N1619;
  assign N1845 = N1835;
  assign N185 = N156;
  assign N211 = N543;
  assign N97 = N1117;
  assign N946 = N48;
  assign N134 = N48;
  assign N1370 = N1536;
  assign N453 = N1536;
  assign N575 = N1536;
  assign N890 = N397;
  assign N613 = N397;
  assign N1021 = N1579;
  assign N737 = N1579;
  assign N741 = N297;
  assign N142 = N297;
  assign N929 = N1466;
  assign N474 = N33;
  assign N1476 = N33;
  assign N1455 = N1794;
  assign N1173 = N146;
  assign N313 = N984;
  assign N284 = N753;
  assign N1062 = N1164;
  assign N39 = N1836;

  CKND2D0BWPHVT U473 ( .A1(N595), .A2(N1203), .ZN(N962) );
  CKND2D0BWPHVT U474 ( .A1(N70), .A2(N505), .ZN(N915) );
  CKND2D0BWPHVT U475 ( .A1(N750), .A2(N506), .ZN(N837) );
  CKND2D0BWPHVT U476 ( .A1(N258), .A2(N227), .ZN(N790) );
  CKND2D0BWPHVT U477 ( .A1(N663), .A2(N249), .ZN(N78) );
  CKND2D0BWPHVT U478 ( .A1(N1352), .A2(N513), .ZN(N750) );
  CKND2D0BWPHVT U479 ( .A1(N1803), .A2(N187), .ZN(N730) );
  CKND2D0BWPHVT U480 ( .A1(N456), .A2(N648), .ZN(N707) );
  AN2D0BWPHVT U481 ( .A1(N442), .A2(N198), .Z(N701) );
  AN2D0BWPHVT U482 ( .A1(N442), .A2(N886), .Z(N700) );
  CKND2D0BWPHVT U483 ( .A1(N1853), .A2(N1181), .ZN(N886) );
  CKND2D0BWPHVT U484 ( .A1(N673), .A2(N287), .ZN(N70) );
  CKND2D0BWPHVT U485 ( .A1(N1343), .A2(N640), .ZN(N676) );
  CKND2D0BWPHVT U486 ( .A1(N769), .A2(N918), .ZN(N664) );
  CKND2D0BWPHVT U487 ( .A1(N786), .A2(N1670), .ZN(N633) );
  CKND2D0BWPHVT U488 ( .A1(N1339), .A2(N1619), .ZN(N618) );
  CKND2D0BWPHVT U489 ( .A1(N677), .A2(N1226), .ZN(N595) );
  CKND2D0BWPHVT U490 ( .A1(N1626), .A2(N1010), .ZN(N558) );
  CKND2D0BWPHVT U491 ( .A1(N171), .A2(N218), .ZN(N555) );
  CKND2D0BWPHVT U492 ( .A1(N94), .A2(N1849), .ZN(N547) );
  CKND2D0BWPHVT U493 ( .A1(N1101), .A2(N1332), .ZN(N94) );
  CKND2D0BWPHVT U494 ( .A1(N842), .A2(N1818), .ZN(N521) );
  CKND2D0BWPHVT U495 ( .A1(N1710), .A2(N340), .ZN(N842) );
  CKND2D0BWPHVT U496 ( .A1(N829), .A2(N868), .ZN(N506) );
  CKND0BWPHVT U497 ( .I(N1352), .ZN(N829) );
  CKND2D0BWPHVT U498 ( .A1(N887), .A2(N218), .ZN(N505) );
  CKND2D0BWPHVT U499 ( .A1(N74), .A2(N36), .ZN(N485) );
  CKND2D0BWPHVT U500 ( .A1(N298), .A2(N124), .ZN(N74) );
  CKND2D0BWPHVT U501 ( .A1(N299), .A2(N909), .ZN(N465) );
  CKND2D0BWPHVT U502 ( .A1(N1708), .A2(N1697), .ZN(N455) );
  AN2D0BWPHVT U503 ( .A1(N442), .A2(N956), .Z(N443) );
  CKND2D0BWPHVT U504 ( .A1(N772), .A2(N1277), .ZN(N956) );
  CKND2D0BWPHVT U505 ( .A1(N1677), .A2(N1107), .ZN(N772) );
  CKND2D0BWPHVT U506 ( .A1(N1674), .A2(N1055), .ZN(N422) );
  CKND2D0BWPHVT U507 ( .A1(N1559), .A2(N108), .ZN(N361) );
  CKND2D0BWPHVT U508 ( .A1(N604), .A2(N21), .ZN(N36) );
  CKND2D0BWPHVT U509 ( .A1(N125), .A2(N2), .ZN(N356) );
  CKND2D0BWPHVT U510 ( .A1(N781), .A2(N1034), .ZN(N346) );
  CKND2D0BWPHVT U511 ( .A1(N95), .A2(N1236), .ZN(N781) );
  CKND2D0BWPHVT U512 ( .A1(N1432), .A2(N651), .ZN(N303) );
  CKND0BWPHVT U513 ( .I(N691), .ZN(N651) );
  CKND2D0BWPHVT U514 ( .A1(N174), .A2(N287), .ZN(N296) );
  CKND2D0BWPHVT U515 ( .A1(N1043), .A2(N528), .ZN(N278) );
  CKND2D0BWPHVT U516 ( .A1(N1000), .A2(N959), .ZN(N25) );
  CKND2D0BWPHVT U517 ( .A1(N416), .A2(N1583), .ZN(N246) );
  CKND2D0BWPHVT U518 ( .A1(N1317), .A2(N945), .ZN(N235) );
  CKND2D0BWPHVT U519 ( .A1(N1765), .A2(N131), .ZN(N230) );
  CKND2D0BWPHVT U520 ( .A1(N1492), .A2(N1488), .ZN(N217) );
  CKND2D0BWPHVT U521 ( .A1(N1817), .A2(N149), .ZN(N198) );
  CKND2D0BWPHVT U522 ( .A1(N809), .A2(N1374), .ZN(N190) );
  CKND2D0BWPHVT U523 ( .A1(N110), .A2(N684), .ZN(N809) );
  CKND2D0BWPHVT U524 ( .A1(N365), .A2(N509), .ZN(N1862) );
  CKND2D0BWPHVT U525 ( .A1(N359), .A2(N947), .ZN(N1853) );
  CKND2D0BWPHVT U526 ( .A1(N1784), .A2(N75), .ZN(N1849) );
  CKND2D0BWPHVT U527 ( .A1(N242), .A2(N1091), .ZN(N1818) );
  CKND2D0BWPHVT U528 ( .A1(N1439), .A2(N1274), .ZN(N1817) );
  CKND2D0BWPHVT U529 ( .A1(N436), .A2(N342), .ZN(N181) );
  AN2D0BWPHVT U530 ( .A1(N442), .A2(N355), .Z(N1804) );
  CKND2D0BWPHVT U531 ( .A1(N85), .A2(N1715), .ZN(N355) );
  CKND2D0BWPHVT U532 ( .A1(N1821), .A2(N1613), .ZN(N85) );
  CKND0BWPHVT U533 ( .I(N1101), .ZN(N1784) );
  CKND2D0BWPHVT U534 ( .A1(N1608), .A2(N29), .ZN(N1765) );
  CKND2D0BWPHVT U535 ( .A1(N862), .A2(N1724), .ZN(N1735) );
  CKND2D0BWPHVT U536 ( .A1(N830), .A2(N1646), .ZN(N862) );
  CKND0BWPHVT U537 ( .I(N1045), .ZN(N830) );
  CKND2D0BWPHVT U538 ( .A1(N162), .A2(N1045), .ZN(N1724) );
  CKND2D0BWPHVT U539 ( .A1(N1180), .A2(N1790), .ZN(N1715) );
  CKND0BWPHVT U540 ( .I(N1821), .ZN(N1790) );
  CKND2D0BWPHVT U541 ( .A1(n419), .A2(N749), .ZN(N1821) );
  CKND2D0BWPHVT U542 ( .A1(N1189), .A2(N227), .ZN(N1708) );
  AN2D0BWPHVT U543 ( .A1(N442), .A2(N1366), .Z(N1703) );
  CKND2D0BWPHVT U544 ( .A1(N1686), .A2(N648), .ZN(N1697) );
  CKND0BWPHVT U545 ( .I(N1189), .ZN(N1686) );
  CKND2D0BWPHVT U546 ( .A1(N996), .A2(N187), .ZN(N1674) );
  CKND2D0BWPHVT U547 ( .A1(N1031), .A2(N1136), .ZN(N1655) );
  CKND0BWPHVT U548 ( .I(N162), .ZN(N1646) );
  CKND2D0BWPHVT U549 ( .A1(N1444), .A2(N1405), .ZN(N1626) );
  CKND2D0BWPHVT U550 ( .A1(N841), .A2(N1527), .ZN(N1620) );
  CKND2D0BWPHVT U551 ( .A1(N1705), .A2(N1502), .ZN(N162) );
  CKND2D0BWPHVT U552 ( .A1(N1141), .A2(N904), .ZN(N1705) );
  CKND2D0BWPHVT U553 ( .A1(N589), .A2(N330), .ZN(N1586) );
  CKND2D0BWPHVT U554 ( .A1(N1168), .A2(N1104), .ZN(N330) );
  CKND2D0BWPHVT U555 ( .A1(N845), .A2(N151), .ZN(N589) );
  CKND0BWPHVT U556 ( .I(N1168), .ZN(N845) );
  CKND2D0BWPHVT U557 ( .A1(N718), .A2(N597), .ZN(N1542) );
  CKND2D0BWPHVT U558 ( .A1(N1625), .A2(N1343), .ZN(N597) );
  CKND2D0BWPHVT U559 ( .A1(N736), .A2(N1074), .ZN(N718) );
  NR2D0BWPHVT U560 ( .A1(N747), .A2(N1630), .ZN(N1515) );
  INR3D0BWPHVT U561 ( .A1(N1011), .B1(N1502), .B2(N77), .ZN(N1630) );
  AN4D0BWPHVT U562 ( .A1(N43), .A2(N1011), .A3(N77), .A4(N428), .Z(N747) );
  INR2D0BWPHVT U563 ( .A1(N1750), .B1(N689), .ZN(N43) );
  AN4D0BWPHVT U564 ( .A1(N1809), .A2(N58), .A3(n420), .A4(n421), .Z(N1750) );
  AN4D0BWPHVT U565 ( .A1(N172), .A2(N1580), .A3(N1280), .A4(N119), .Z(n421) );
  ND3D0BWPHVT U566 ( .A1(n422), .A2(N1490), .A3(N489), .ZN(N1580) );
  NR2D0BWPHVT U567 ( .A1(N1130), .A2(N1360), .ZN(N489) );
  ND3D0BWPHVT U568 ( .A1(N1490), .A2(N1802), .A3(n422), .ZN(N172) );
  AN2D0BWPHVT U569 ( .A1(N832), .A2(N606), .Z(n420) );
  ND3D0BWPHVT U570 ( .A1(N1727), .A2(N175), .A3(n422), .ZN(N606) );
  ND3D0BWPHVT U571 ( .A1(N1054), .A2(N1294), .A3(n423), .ZN(N832) );
  ND3D0BWPHVT U572 ( .A1(N1054), .A2(N495), .A3(n423), .ZN(N58) );
  ND3D0BWPHVT U573 ( .A1(n423), .A2(N1124), .A3(N856), .ZN(N1809) );
  NR2D0BWPHVT U574 ( .A1(N1645), .A2(N543), .ZN(N856) );
  CKND2D0BWPHVT U575 ( .A1(N1252), .A2(N1521), .ZN(N1500) );
  CKND2D0BWPHVT U576 ( .A1(N898), .A2(N528), .ZN(N1492) );
  CKND2D0BWPHVT U577 ( .A1(N1394), .A2(N752), .ZN(N149) );
  CKND0BWPHVT U578 ( .I(N1274), .ZN(N752) );
  CKND2D0BWPHVT U579 ( .A1(N734), .A2(N338), .ZN(N1488) );
  CKND2D0BWPHVT U580 ( .A1(N1525), .A2(N1369), .ZN(N1459) );
  AN2D0BWPHVT U581 ( .A1(N442), .A2(N725), .Z(N1442) );
  CKND2D0BWPHVT U582 ( .A1(N306), .A2(N1510), .ZN(N725) );
  CKND2D0BWPHVT U583 ( .A1(N1658), .A2(N1233), .ZN(N1510) );
  CKND2D0BWPHVT U584 ( .A1(N1269), .A2(N1234), .ZN(N306) );
  CKND2D0BWPHVT U585 ( .A1(N1502), .A2(N127), .ZN(N442) );
  CKND2D0BWPHVT U586 ( .A1(N458), .A2(N124), .ZN(N1434) );
  CKND2D0BWPHVT U587 ( .A1(N1252), .A2(N1307), .ZN(N1415) );
  CKND2D0BWPHVT U588 ( .A1(N526), .A2(N1414), .ZN(N1396) );
  CKND2D0BWPHVT U589 ( .A1(N884), .A2(N1706), .ZN(N1390) );
  CKND2D0BWPHVT U590 ( .A1(N273), .A2(N1000), .ZN(N1706) );
  CKND2D0BWPHVT U591 ( .A1(N153), .A2(N416), .ZN(N884) );
  CKND2D0BWPHVT U592 ( .A1(N1307), .A2(N316), .ZN(N1389) );
  CKND2D0BWPHVT U593 ( .A1(N1297), .A2(N588), .ZN(N138) );
  CKND2D0BWPHVT U594 ( .A1(N977), .A2(N876), .ZN(N1374) );
  CKND2D0BWPHVT U595 ( .A1(N889), .A2(N1129), .ZN(N1366) );
  CKND2D0BWPHVT U596 ( .A1(N440), .A2(N1327), .ZN(N889) );
  CKND2D0BWPHVT U597 ( .A1(N225), .A2(N338), .ZN(N1341) );
  CKND2D0BWPHVT U598 ( .A1(N1074), .A2(N49), .ZN(N1337) );
  CKND2D0BWPHVT U599 ( .A1(N1422), .A2(N1136), .ZN(N131) );
  ND3D0BWPHVT U600 ( .A1(N1124), .A2(N374), .A3(n423), .ZN(N1280) );
  AN3D0BWPHVT U601 ( .A1(N1490), .A2(N270), .A3(N1727), .Z(n423) );
  CKND2D0BWPHVT U602 ( .A1(N1612), .A2(N1383), .ZN(N1277) );
  CKND0BWPHVT U603 ( .I(N1677), .ZN(N1383) );
  CKND0BWPHVT U604 ( .I(N1107), .ZN(N1612) );
  CKND2D0BWPHVT U605 ( .A1(n419), .A2(N949), .ZN(N1274) );
  CKND0BWPHVT U606 ( .I(N77), .ZN(N127) );
  CKND2D0BWPHVT U607 ( .A1(N352), .A2(N1663), .ZN(N1263) );
  CKND2D0BWPHVT U608 ( .A1(N1588), .A2(N2), .ZN(N1663) );
  CKND2D0BWPHVT U609 ( .A1(N1795), .A2(N509), .ZN(N352) );
  CKND2D0BWPHVT U610 ( .A1(N231), .A2(N1236), .ZN(N1253) );
  CKND0BWPHVT U611 ( .I(N1233), .ZN(N1234) );
  CKND2D0BWPHVT U612 ( .A1(n419), .A2(N1265), .ZN(N1233) );
  CKND2D0BWPHVT U613 ( .A1(N805), .A2(N311), .ZN(N121) );
  CKND2D0BWPHVT U614 ( .A1(N1828), .A2(N1317), .ZN(N1207) );
  CKND2D0BWPHVT U615 ( .A1(N1570), .A2(N429), .ZN(N1203) );
  CKND0BWPHVT U616 ( .I(N677), .ZN(N429) );
  CKND2D0BWPHVT U617 ( .A1(N791), .A2(N1502), .ZN(N677) );
  CKND2D0BWPHVT U618 ( .A1(N1053), .A2(N1048), .ZN(N791) );
  CKND0BWPHVT U619 ( .I(N1226), .ZN(N1570) );
  CKND2D0BWPHVT U620 ( .A1(N680), .A2(N1610), .ZN(N1226) );
  CKND2D0BWPHVT U621 ( .A1(N1026), .A2(N1223), .ZN(N1610) );
  CKND2D0BWPHVT U622 ( .A1(N32), .A2(N632), .ZN(N680) );
  CKND0BWPHVT U623 ( .I(N1223), .ZN(N632) );
  CKND2D0BWPHVT U624 ( .A1(N1598), .A2(N1369), .ZN(N1223) );
  ND3D0BWPHVT U625 ( .A1(N1727), .A2(N539), .A3(n422), .ZN(N119) );
  AN3D0BWPHVT U626 ( .A1(N1124), .A2(N270), .A3(N1054), .Z(n422) );
  CKND0BWPHVT U627 ( .I(N106), .ZN(N270) );
  CKND2D0BWPHVT U628 ( .A1(N206), .A2(N21), .ZN(N1185) );
  CKND2D0BWPHVT U629 ( .A1(N1097), .A2(N945), .ZN(N1183) );
  CKND2D0BWPHVT U630 ( .A1(N1354), .A2(N1356), .ZN(N1181) );
  CKND0BWPHVT U631 ( .I(N359), .ZN(N1354) );
  XNR2D0BWPHVT U632 ( .A1(N588), .A2(N1297), .ZN(N359) );
  CKND0BWPHVT U633 ( .I(N311), .ZN(N588) );
  CKND2D0BWPHVT U634 ( .A1(n419), .A2(N882), .ZN(N311) );
  CKND0BWPHVT U635 ( .I(N1613), .ZN(N1180) );
  CKND2D0BWPHVT U636 ( .A1(N814), .A2(N1367), .ZN(N1129) );
  CKND0BWPHVT U637 ( .I(N440), .ZN(N1367) );
  CKND0BWPHVT U638 ( .I(N1327), .ZN(N814) );
  CKND2D0BWPHVT U639 ( .A1(n419), .A2(N678), .ZN(N1327) );
  CKND2D0BWPHVT U640 ( .A1(N608), .A2(N29), .ZN(N1115) );
  CKND2D0BWPHVT U641 ( .A1(n419), .A2(N502), .ZN(N1107) );
  NR2D0BWPHVT U642 ( .A1(n424), .A2(N480), .ZN(n419) );
  CKND0BWPHVT U643 ( .I(N689), .ZN(n424) );
  CKND2D0BWPHVT U644 ( .A1(N350), .A2(N666), .ZN(N689) );
  CKND0BWPHVT U645 ( .I(N20), .ZN(N666) );
  CKND0BWPHVT U646 ( .I(N1296), .ZN(N350) );
  CKND2D0BWPHVT U647 ( .A1(N704), .A2(N691), .ZN(N11) );
  CKND0BWPHVT U648 ( .I(N1828), .ZN(N108) );
  CKND2D0BWPHVT U649 ( .A1(N1213), .A2(N249), .ZN(N1055) );
  CKND2D0BWPHVT U650 ( .A1(N1559), .A2(N1521), .ZN(N1046) );
  CKND2D0BWPHVT U651 ( .A1(N1852), .A2(N1002), .ZN(N1045) );
  CKND2D0BWPHVT U652 ( .A1(N1448), .A2(N503), .ZN(N1852) );
  CKND0BWPHVT U653 ( .I(N1190), .ZN(N1448) );
  CKND2D0BWPHVT U654 ( .A1(N973), .A2(N1670), .ZN(N1034) );
  CKND0BWPHVT U655 ( .I(N32), .ZN(N1026) );
  CKND2D0BWPHVT U656 ( .A1(N428), .A2(N20), .ZN(N32) );
  ND4D0BWPHVT U657 ( .A1(N1168), .A2(N1352), .A3(n425), .A4(n426), .ZN(N20) );
  NR4D0BWPHVT U658 ( .A1(N996), .A2(N887), .A3(N604), .A4(N1795), .ZN(n426) );
  CKND0BWPHVT U659 ( .I(N1588), .ZN(N1795) );
  ND3D0BWPHVT U660 ( .A1(N495), .A2(n427), .A3(N1490), .ZN(N1588) );
  CKND0BWPHVT U661 ( .I(N298), .ZN(N604) );
  ND3D0BWPHVT U662 ( .A1(N1294), .A2(N539), .A3(n428), .ZN(N298) );
  CKND0BWPHVT U663 ( .I(N673), .ZN(N887) );
  ND3D0BWPHVT U664 ( .A1(N1294), .A2(n427), .A3(N1490), .ZN(N673) );
  CKND0BWPHVT U665 ( .I(N1213), .ZN(N996) );
  ND3D0BWPHVT U666 ( .A1(N1124), .A2(n427), .A3(N539), .ZN(N1213) );
  NR2D0BWPHVT U667 ( .A1(N1114), .A2(N1608), .ZN(n425) );
  CKND0BWPHVT U668 ( .I(N1422), .ZN(N1608) );
  ND3D0BWPHVT U669 ( .A1(N1124), .A2(n427), .A3(N175), .ZN(N1422) );
  AN3D0BWPHVT U670 ( .A1(N1802), .A2(N600), .A3(N374), .Z(n427) );
  ND3D0BWPHVT U671 ( .A1(N495), .A2(N539), .A3(n428), .ZN(N1352) );
  ND3D0BWPHVT U672 ( .A1(n428), .A2(N1490), .A3(N1493), .ZN(N1168) );
  ND4D0BWPHVT U673 ( .A1(N1727), .A2(N1054), .A3(N1490), .A4(N1124), .ZN(N1011) );
  NR2D0BWPHVT U674 ( .A1(N1861), .A2(N581), .ZN(N1490) );
  CKND2D0BWPHVT U675 ( .A1(N1114), .A2(N1073), .ZN(N1010) );
  CKND0BWPHVT U676 ( .I(N1444), .ZN(N1114) );
  ND3D0BWPHVT U677 ( .A1(N66), .A2(N1124), .A3(n428), .ZN(N1444) );
  AN3D0BWPHVT U678 ( .A1(N1802), .A2(N600), .A3(N1054), .Z(n428) );
  CKND2D0BWPHVT U679 ( .A1(N789), .A2(N106), .ZN(N600) );
  ND3D0BWPHVT U680 ( .A1(n429), .A2(N1273), .A3(N437), .ZN(N789) );
  CKND0BWPHVT U681 ( .I(N1598), .ZN(n429) );
  CKND2D0BWPHVT U682 ( .A1(N1502), .A2(N519), .ZN(N1598) );
  CKND0BWPHVT U683 ( .I(N1048), .ZN(N519) );
  CKND2D0BWPHVT U684 ( .A1(N909), .A2(N1097), .ZN(N1009) );
  CKND2D0BWPHVT U685 ( .A1(N1190), .A2(N568), .ZN(N1002) );
  CKND0BWPHVT U686 ( .I(N503), .ZN(N568) );
  CKND2D0BWPHVT U687 ( .A1(N780), .A2(N176), .ZN(N503) );
  CKND0BWPHVT U688 ( .I(N305), .ZN(N176) );
  CKND2D0BWPHVT U689 ( .A1(N38), .A2(N1632), .ZN(N305) );
  CKND2D0BWPHVT U690 ( .A1(N299), .A2(N290), .ZN(N1632) );
  CKND2D0BWPHVT U691 ( .A1(N316), .A2(N1536), .ZN(N38) );
  CKND0BWPHVT U692 ( .I(N299), .ZN(N316) );
  CKND2D0BWPHVT U693 ( .A1(N1296), .A2(N428), .ZN(N1190) );
  ND4D0BWPHVT U694 ( .A1(N1101), .A2(N1189), .A3(n430), .A4(n431), .ZN(N1296)
         );
  NR4D0BWPHVT U695 ( .A1(N977), .A2(N95), .A3(N734), .A4(N1625), .ZN(n431) );
  CKND0BWPHVT U696 ( .I(N736), .ZN(N1625) );
  ND3D0BWPHVT U697 ( .A1(N66), .A2(N1124), .A3(n432), .ZN(N736) );
  NR2D0BWPHVT U698 ( .A1(N1), .A2(N1589), .ZN(N1124) );
  CKND0BWPHVT U699 ( .I(N898), .ZN(N734) );
  ND3D0BWPHVT U700 ( .A1(N495), .A2(N539), .A3(n432), .ZN(N898) );
  CKND0BWPHVT U701 ( .I(N973), .ZN(N95) );
  ND3D0BWPHVT U702 ( .A1(N66), .A2(n433), .A3(N495), .ZN(N973) );
  NR2D0BWPHVT U703 ( .A1(N1324), .A2(N1589), .ZN(N495) );
  CKND0BWPHVT U704 ( .I(N110), .ZN(N977) );
  ND3D0BWPHVT U705 ( .A1(N1294), .A2(n433), .A3(N66), .ZN(N110) );
  NR2D0BWPHVT U706 ( .A1(N928), .A2(N368), .ZN(N66) );
  NR2D0BWPHVT U707 ( .A1(N1710), .A2(N273), .ZN(n430) );
  CKND0BWPHVT U708 ( .I(N153), .ZN(N273) );
  ND3D0BWPHVT U709 ( .A1(n433), .A2(N539), .A3(N1493), .ZN(N153) );
  NR2D0BWPHVT U710 ( .A1(N1324), .A2(N30), .ZN(N1493) );
  CKND0BWPHVT U711 ( .I(N1), .ZN(N1324) );
  AN3D0BWPHVT U712 ( .A1(N1802), .A2(N10), .A3(N374), .Z(n433) );
  CKND0BWPHVT U713 ( .I(N242), .ZN(N1710) );
  ND4D0BWPHVT U714 ( .A1(N1802), .A2(N10), .A3(N1294), .A4(n434), .ZN(N242) );
  AN2D0BWPHVT U715 ( .A1(N1054), .A2(N175), .Z(n434) );
  NR2D0BWPHVT U716 ( .A1(N1820), .A2(N1645), .ZN(N1054) );
  NR2D0BWPHVT U717 ( .A1(N709), .A2(N240), .ZN(N1802) );
  CKND0BWPHVT U718 ( .I(N1360), .ZN(N240) );
  ND3D0BWPHVT U719 ( .A1(N1294), .A2(N539), .A3(n432), .ZN(N1189) );
  NR2D0BWPHVT U720 ( .A1(N368), .A2(N1861), .ZN(N539) );
  CKND0BWPHVT U721 ( .I(N581), .ZN(N368) );
  ND3D0BWPHVT U722 ( .A1(N175), .A2(N1294), .A3(n432), .ZN(N1101) );
  AN3D0BWPHVT U723 ( .A1(N374), .A2(N10), .A3(N1727), .Z(n432) );
  NR2D0BWPHVT U724 ( .A1(N709), .A2(N1360), .ZN(N1727) );
  CKND2D0BWPHVT U725 ( .A1(N1729), .A2(N1221), .ZN(N1360) );
  CKND2D0BWPHVT U726 ( .A1(N502), .A2(N1783), .ZN(N1221) );
  CKND0BWPHVT U727 ( .I(N297), .ZN(N502) );
  CKND2D0BWPHVT U728 ( .A1(N297), .A2(N1801), .ZN(N1729) );
  CKND0BWPHVT U729 ( .I(N1783), .ZN(N1801) );
  CKND2D0BWPHVT U730 ( .A1(N1677), .A2(N480), .ZN(N1783) );
  CKND2D0BWPHVT U731 ( .A1(N636), .A2(N1713), .ZN(N1677) );
  CKND2D0BWPHVT U732 ( .A1(N1527), .A2(N1369), .ZN(N1713) );
  CKND0BWPHVT U733 ( .I(N841), .ZN(N1369) );
  CKND2D0BWPHVT U734 ( .A1(N841), .A2(N1525), .ZN(N636) );
  CKND0BWPHVT U735 ( .I(N1527), .ZN(N1525) );
  CKND2D0BWPHVT U736 ( .A1(N239), .A2(N1039), .ZN(N1527) );
  CKND2D0BWPHVT U737 ( .A1(N1604), .A2(N1078), .ZN(N1039) );
  CKND0BWPHVT U738 ( .I(N1298), .ZN(N1078) );
  CKND0BWPHVT U739 ( .I(N1117), .ZN(N1604) );
  CKND2D0BWPHVT U740 ( .A1(N1298), .A2(N1117), .ZN(N239) );
  CKND2D0BWPHVT U741 ( .A1(N1053), .A2(N428), .ZN(N1117) );
  CKND2D0BWPHVT U742 ( .A1(N907), .A2(N1462), .ZN(N1298) );
  CKND2D0BWPHVT U743 ( .A1(N1521), .A2(N1091), .ZN(N1462) );
  CKND2D0BWPHVT U744 ( .A1(N945), .A2(N340), .ZN(N907) );
  CKND0BWPHVT U745 ( .I(N1521), .ZN(N945) );
  CKND2D0BWPHVT U746 ( .A1(N1591), .A2(N1393), .ZN(N841) );
  CKND2D0BWPHVT U747 ( .A1(N309), .A2(N490), .ZN(N1393) );
  CKND0BWPHVT U748 ( .I(N1579), .ZN(N490) );
  CKND2D0BWPHVT U749 ( .A1(N1139), .A2(N1579), .ZN(N1591) );
  CKND2D0BWPHVT U750 ( .A1(N788), .A2(N1428), .ZN(N1579) );
  CKND2D0BWPHVT U751 ( .A1(N1104), .A2(N29), .ZN(N1428) );
  CKND2D0BWPHVT U752 ( .A1(N1136), .A2(N151), .ZN(N788) );
  CKND0BWPHVT U753 ( .I(N309), .ZN(N1139) );
  XNR2D0BWPHVT U754 ( .A1(N1252), .A2(N909), .ZN(N309) );
  CKND2D0BWPHVT U755 ( .A1(N1126), .A2(N683), .ZN(N297) );
  CKND0BWPHVT U756 ( .I(N1130), .ZN(N709) );
  CKND2D0BWPHVT U757 ( .A1(N241), .A2(N683), .ZN(N1130) );
  CKND2D0BWPHVT U758 ( .A1(N708), .A2(N480), .ZN(N683) );
  NR2D0BWPHVT U759 ( .A1(N357), .A2(N1820), .ZN(N374) );
  CKND0BWPHVT U760 ( .I(N543), .ZN(N1820) );
  CKND2D0BWPHVT U761 ( .A1(N767), .A2(N427), .ZN(N543) );
  CKND0BWPHVT U762 ( .I(N1645), .ZN(N357) );
  CKND2D0BWPHVT U763 ( .A1(N1709), .A2(N1692), .ZN(N1645) );
  CKND2D0BWPHVT U764 ( .A1(N638), .A2(N1449), .ZN(N1692) );
  CKND0BWPHVT U765 ( .I(N749), .ZN(N1449) );
  CKND0BWPHVT U766 ( .I(N1018), .ZN(N638) );
  CKND2D0BWPHVT U767 ( .A1(N749), .A2(N1018), .ZN(N1709) );
  CKND2D0BWPHVT U768 ( .A1(N1613), .A2(N480), .ZN(N1018) );
  CKND2D0BWPHVT U769 ( .A1(N966), .A2(N825), .ZN(N1613) );
  CKND2D0BWPHVT U770 ( .A1(N628), .A2(N33), .ZN(N825) );
  CKND2D0BWPHVT U771 ( .A1(N1760), .A2(N745), .ZN(N966) );
  CKND0BWPHVT U772 ( .I(N33), .ZN(N745) );
  CKND2D0BWPHVT U773 ( .A1(N1794), .A2(N146), .ZN(N33) );
  CKND2D0BWPHVT U774 ( .A1(N1035), .A2(N779), .ZN(N146) );
  CKND0BWPHVT U775 ( .I(N984), .ZN(N779) );
  CKND0BWPHVT U776 ( .I(N1836), .ZN(N1035) );
  CKND2D0BWPHVT U777 ( .A1(N984), .A2(N1836), .ZN(N1794) );
  CKND2D0BWPHVT U778 ( .A1(N1141), .A2(N428), .ZN(N1836) );
  CKND2D0BWPHVT U779 ( .A1(N753), .A2(N1164), .ZN(N984) );
  CKND2D0BWPHVT U780 ( .A1(N1332), .A2(N29), .ZN(N1164) );
  CKND2D0BWPHVT U781 ( .A1(N1136), .A2(N75), .ZN(N753) );
  CKND0BWPHVT U782 ( .I(N628), .ZN(N1760) );
  XNR2D0BWPHVT U783 ( .A1(N1828), .A2(N1317), .ZN(N628) );
  XNR2D0BWPHVT U784 ( .A1(N1521), .A2(N1097), .ZN(N1828) );
  CKND0BWPHVT U785 ( .I(N1252), .ZN(N1097) );
  XNR2D0BWPHVT U786 ( .A1(N1803), .A2(N187), .ZN(N1252) );
  CKND0BWPHVT U787 ( .I(N663), .ZN(N1803) );
  CKND2D0BWPHVT U788 ( .A1(N687), .A2(N1700), .ZN(N663) );
  CKND2D0BWPHVT U789 ( .A1(N287), .A2(N509), .ZN(N1700) );
  CKND2D0BWPHVT U790 ( .A1(N2), .A2(N218), .ZN(N687) );
  NR2D0BWPHVT U791 ( .A1(N30), .A2(N1), .ZN(N1294) );
  CKND0BWPHVT U792 ( .I(N1589), .ZN(N30) );
  CKND2D0BWPHVT U793 ( .A1(N1261), .A2(N1162), .ZN(N1589) );
  CKND2D0BWPHVT U794 ( .A1(N112), .A2(N590), .ZN(N1162) );
  CKND0BWPHVT U795 ( .I(N949), .ZN(N590) );
  CKND0BWPHVT U796 ( .I(N1806), .ZN(N112) );
  CKND2D0BWPHVT U797 ( .A1(N1806), .A2(N949), .ZN(N1261) );
  CKND2D0BWPHVT U798 ( .A1(N1439), .A2(N480), .ZN(N1806) );
  CKND0BWPHVT U799 ( .I(N1394), .ZN(N1439) );
  XNR2D0BWPHVT U800 ( .A1(N342), .A2(N769), .ZN(N1394) );
  CKND0BWPHVT U801 ( .I(N436), .ZN(N769) );
  XNR2D0BWPHVT U802 ( .A1(N171), .A2(N218), .ZN(N436) );
  CKND0BWPHVT U803 ( .I(N287), .ZN(N218) );
  CKND0BWPHVT U804 ( .I(N174), .ZN(N171) );
  CKND2D0BWPHVT U805 ( .A1(N751), .A2(N1007), .ZN(N174) );
  CKND2D0BWPHVT U806 ( .A1(N124), .A2(N151), .ZN(N1007) );
  CKND2D0BWPHVT U807 ( .A1(N1104), .A2(N21), .ZN(N751) );
  CKND0BWPHVT U808 ( .I(N918), .ZN(N342) );
  CKND2D0BWPHVT U809 ( .A1(N1446), .A2(N1085), .ZN(N918) );
  CKND2D0BWPHVT U810 ( .A1(N697), .A2(N1414), .ZN(N1085) );
  CKND2D0BWPHVT U811 ( .A1(N1619), .A2(N329), .ZN(N1446) );
  CKND0BWPHVT U812 ( .I(N697), .ZN(N329) );
  CKND2D0BWPHVT U813 ( .A1(N461), .A2(N1040), .ZN(N697) );
  CKND2D0BWPHVT U814 ( .A1(N646), .A2(N648), .ZN(N1040) );
  CKND2D0BWPHVT U815 ( .A1(N953), .A2(N227), .ZN(N461) );
  CKND0BWPHVT U816 ( .I(N646), .ZN(N953) );
  XNR2D0BWPHVT U817 ( .A1(N1583), .A2(N1000), .ZN(N646) );
  CKND0BWPHVT U818 ( .I(N959), .ZN(N1583) );
  ND3D0BWPHVT U819 ( .A1(N428), .A2(N708), .A3(N241), .ZN(N959) );
  NR2D0BWPHVT U820 ( .A1(N928), .A2(N581), .ZN(N175) );
  CKND2D0BWPHVT U821 ( .A1(N89), .A2(N1830), .ZN(N581) );
  CKND2D0BWPHVT U822 ( .A1(N93), .A2(N1693), .ZN(N1830) );
  CKND0BWPHVT U823 ( .I(N882), .ZN(N1693) );
  CKND0BWPHVT U824 ( .I(N596), .ZN(N93) );
  CKND2D0BWPHVT U825 ( .A1(N596), .A2(N882), .ZN(N89) );
  CKND2D0BWPHVT U826 ( .A1(N480), .A2(N1119), .ZN(N596) );
  CKND2D0BWPHVT U827 ( .A1(N1413), .A2(N1125), .ZN(N1119) );
  CKND2D0BWPHVT U828 ( .A1(N805), .A2(N947), .ZN(N1125) );
  CKND0BWPHVT U829 ( .I(N1356), .ZN(N947) );
  CKND2D0BWPHVT U830 ( .A1(N1297), .A2(N1356), .ZN(N1413) );
  CKND2D0BWPHVT U831 ( .A1(N1541), .A2(N1437), .ZN(N1356) );
  CKND2D0BWPHVT U832 ( .A1(N1840), .A2(N249), .ZN(N1437) );
  CKND0BWPHVT U833 ( .I(N1466), .ZN(N1840) );
  CKND2D0BWPHVT U834 ( .A1(N187), .A2(N1466), .ZN(N1541) );
  ND3D0BWPHVT U835 ( .A1(N428), .A2(N708), .A3(N1126), .ZN(N1466) );
  CKND0BWPHVT U836 ( .I(N1653), .ZN(N708) );
  CKND0BWPHVT U837 ( .I(N249), .ZN(N187) );
  CKND0BWPHVT U838 ( .I(N805), .ZN(N1297) );
  XNR2D0BWPHVT U839 ( .A1(N299), .A2(N909), .ZN(N805) );
  CKND0BWPHVT U840 ( .I(N1307), .ZN(N909) );
  XNR2D0BWPHVT U841 ( .A1(N206), .A2(N21), .ZN(N1307) );
  CKND0BWPHVT U842 ( .I(N124), .ZN(N21) );
  CKND0BWPHVT U843 ( .I(N458), .ZN(N206) );
  CKND2D0BWPHVT U844 ( .A1(N1834), .A2(N1245), .ZN(N458) );
  CKND2D0BWPHVT U845 ( .A1(N513), .A2(N1073), .ZN(N1245) );
  CKND2D0BWPHVT U846 ( .A1(N1405), .A2(N868), .ZN(N1834) );
  XNR2D0BWPHVT U847 ( .A1(N1521), .A2(N1317), .ZN(N299) );
  CKND0BWPHVT U848 ( .I(N1559), .ZN(N1317) );
  XNR2D0BWPHVT U849 ( .A1(N456), .A2(N648), .ZN(N1559) );
  CKND0BWPHVT U850 ( .I(N227), .ZN(N648) );
  CKND0BWPHVT U851 ( .I(N258), .ZN(N456) );
  CKND2D0BWPHVT U852 ( .A1(N974), .A2(N727), .ZN(N258) );
  CKND2D0BWPHVT U853 ( .A1(N528), .A2(N1343), .ZN(N727) );
  CKND2D0BWPHVT U854 ( .A1(N1074), .A2(N338), .ZN(N974) );
  XNR2D0BWPHVT U855 ( .A1(N231), .A2(N1236), .ZN(N1521) );
  CKND0BWPHVT U856 ( .I(N786), .ZN(N231) );
  CKND2D0BWPHVT U857 ( .A1(N642), .A2(N1425), .ZN(N786) );
  CKND2D0BWPHVT U858 ( .A1(N684), .A2(N1000), .ZN(N1425) );
  CKND2D0BWPHVT U859 ( .A1(N416), .A2(N876), .ZN(N642) );
  CKND0BWPHVT U860 ( .I(N1861), .ZN(N928) );
  CKND2D0BWPHVT U861 ( .A1(N746), .A2(N661), .ZN(N1861) );
  CKND2D0BWPHVT U862 ( .A1(N1069), .A2(N964), .ZN(N661) );
  CKND0BWPHVT U863 ( .I(N1441), .ZN(N964) );
  CKND2D0BWPHVT U864 ( .A1(N1265), .A2(N1441), .ZN(N746) );
  CKND2D0BWPHVT U865 ( .A1(N1658), .A2(N480), .ZN(N1441) );
  CKND0BWPHVT U866 ( .I(N1269), .ZN(N1658) );
  XNR2D0BWPHVT U867 ( .A1(N691), .A2(N1432), .ZN(N1269) );
  CKND0BWPHVT U868 ( .I(N704), .ZN(N1432) );
  XNR2D0BWPHVT U869 ( .A1(N49), .A2(N1343), .ZN(N704) );
  CKND0BWPHVT U870 ( .I(N1074), .ZN(N1343) );
  CKND0BWPHVT U871 ( .I(N640), .ZN(N49) );
  ND3D0BWPHVT U872 ( .A1(N1134), .A2(N428), .A3(N767), .ZN(N640) );
  XNR2D0BWPHVT U873 ( .A1(N1414), .A2(N1339), .ZN(N691) );
  CKND0BWPHVT U874 ( .I(N526), .ZN(N1339) );
  XNR2D0BWPHVT U875 ( .A1(N608), .A2(N29), .ZN(N526) );
  CKND0BWPHVT U876 ( .I(N1136), .ZN(N29) );
  CKND0BWPHVT U877 ( .I(N1031), .ZN(N608) );
  CKND2D0BWPHVT U878 ( .A1(N798), .A2(N1022), .ZN(N1031) );
  CKND2D0BWPHVT U879 ( .A1(N1670), .A2(N1073), .ZN(N1022) );
  CKND0BWPHVT U880 ( .I(N1405), .ZN(N1073) );
  CKND2D0BWPHVT U881 ( .A1(N1405), .A2(N1236), .ZN(N798) );
  CKND0BWPHVT U882 ( .I(N1619), .ZN(N1414) );
  CKND2D0BWPHVT U883 ( .A1(N1835), .A2(N156), .ZN(N1619) );
  CKND2D0BWPHVT U884 ( .A1(N290), .A2(N876), .ZN(N156) );
  CKND0BWPHVT U885 ( .I(N684), .ZN(N876) );
  CKND0BWPHVT U886 ( .I(N1536), .ZN(N290) );
  CKND2D0BWPHVT U887 ( .A1(N1536), .A2(N684), .ZN(N1835) );
  CKND2D0BWPHVT U888 ( .A1(N48), .A2(N397), .ZN(N1536) );
  CKND2D0BWPHVT U889 ( .A1(N1332), .A2(N340), .ZN(N397) );
  CKND0BWPHVT U890 ( .I(N1091), .ZN(N340) );
  CKND2D0BWPHVT U891 ( .A1(N1091), .A2(N75), .ZN(N48) );
  CKND0BWPHVT U892 ( .I(N1332), .ZN(N75) );
  CKND0BWPHVT U893 ( .I(N1069), .ZN(N1265) );
  CKND2D0BWPHVT U894 ( .A1(N328), .A2(N427), .ZN(N1069) );
  CKND2D0BWPHVT U895 ( .A1(N1134), .A2(N480), .ZN(N427) );
  CKND2D0BWPHVT U896 ( .A1(N905), .A2(N106), .ZN(N10) );
  ND3D0BWPHVT U897 ( .A1(N77), .A2(N428), .A3(N437), .ZN(N106) );
  ND3D0BWPHVT U898 ( .A1(N1273), .A2(n435), .A3(N437), .ZN(N905) );
  CKND2D0BWPHVT U899 ( .A1(N1134), .A2(N1653), .ZN(N437) );
  CKND0BWPHVT U900 ( .I(N780), .ZN(n435) );
  CKND2D0BWPHVT U901 ( .A1(N1502), .A2(N936), .ZN(N780) );
  CKND0BWPHVT U902 ( .I(N904), .ZN(N936) );
  CKND2D0BWPHVT U903 ( .A1(N1745), .A2(N1208), .ZN(N1) );
  CKND2D0BWPHVT U904 ( .A1(N1407), .A2(N1666), .ZN(N1208) );
  CKND0BWPHVT U905 ( .I(N678), .ZN(N1666) );
  CKND0BWPHVT U906 ( .I(N1319), .ZN(N1407) );
  CKND2D0BWPHVT U907 ( .A1(N678), .A2(N1319), .ZN(N1745) );
  CKND2D0BWPHVT U908 ( .A1(N440), .A2(N480), .ZN(N1319) );
  CKND0BWPHVT U909 ( .I(N1273), .ZN(N480) );
  CKND2D0BWPHVT U910 ( .A1(N1160), .A2(N1041), .ZN(N440) );
  CKND2D0BWPHVT U911 ( .A1(N975), .A2(N1637), .ZN(N1041) );
  CKND0BWPHVT U912 ( .I(N504), .ZN(N1637) );
  CKND0BWPHVT U913 ( .I(N1105), .ZN(N975) );
  CKND2D0BWPHVT U914 ( .A1(N504), .A2(N1105), .ZN(N1160) );
  ND3D0BWPHVT U915 ( .A1(N1134), .A2(N428), .A3(N328), .ZN(N1105) );
  CKND0BWPHVT U916 ( .I(N1502), .ZN(N428) );
  CKND2D0BWPHVT U917 ( .A1(N902), .A2(N508), .ZN(N504) );
  CKND2D0BWPHVT U918 ( .A1(N579), .A2(N1505), .ZN(N508) );
  CKND0BWPHVT U919 ( .I(N1196), .ZN(N1505) );
  CKND2D0BWPHVT U920 ( .A1(N1196), .A2(N1123), .ZN(N902) );
  CKND0BWPHVT U921 ( .I(N579), .ZN(N1123) );
  XNR2D0BWPHVT U922 ( .A1(N365), .A2(N509), .ZN(N579) );
  CKND0BWPHVT U923 ( .I(N2), .ZN(N509) );
  CKND0BWPHVT U924 ( .I(N125), .ZN(N365) );
  CKND2D0BWPHVT U925 ( .A1(N872), .A2(N420), .ZN(N125) );
  CKND2D0BWPHVT U926 ( .A1(N513), .A2(N151), .ZN(N420) );
  CKND0BWPHVT U927 ( .I(N1104), .ZN(N151) );
  CKND2D0BWPHVT U928 ( .A1(N1104), .A2(N868), .ZN(N872) );
  CKND0BWPHVT U929 ( .I(N513), .ZN(N868) );
  XNR2D0BWPHVT U930 ( .A1(N225), .A2(N338), .ZN(N1196) );
  CKND0BWPHVT U931 ( .I(N528), .ZN(N338) );
  CKND0BWPHVT U932 ( .I(N1043), .ZN(N225) );
  CKND2D0BWPHVT U933 ( .A1(N388), .A2(N169), .ZN(N1043) );
  CKND2D0BWPHVT U934 ( .A1(N416), .A2(N1236), .ZN(N169) );
  CKND0BWPHVT U935 ( .I(N1670), .ZN(N1236) );
  CKND2D0BWPHVT U936 ( .A1(N1670), .A2(N1000), .ZN(N388) );
  CKND0BWPHVT U937 ( .I(N416), .ZN(N1000) );
endmodule

